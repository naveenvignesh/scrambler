
module se8 ( clk, rst, write, addr, lfsrdin, pushin, datain, entrophy, pushout, 
        dataout );
  input [11:0] addr;
  input [31:0] lfsrdin;
  input [7:0] datain;
  input [31:0] entrophy;
  output [31:0] dataout;
  input clk, rst, write, pushin;
  output pushout;
  wire   \dataselector_shifted[0] , n8684, n8685, n8686, n8687, n8688, n8689,
         n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699,
         n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709,
         n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719,
         n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729,
         n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739,
         n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749,
         n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759,
         n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769,
         n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779,
         n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789,
         n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799,
         n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809,
         n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819,
         n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829,
         n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839,
         n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849,
         n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859,
         n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869,
         n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879,
         n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889,
         n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899,
         n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909,
         n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919,
         n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929,
         n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939,
         n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949,
         n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959,
         n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969,
         n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979,
         n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989,
         n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999,
         n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009,
         n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019,
         n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029,
         n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039,
         n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049,
         n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059,
         n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069,
         n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079,
         n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089,
         n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099,
         n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109,
         n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119,
         n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129,
         n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139,
         n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149,
         n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159,
         n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169,
         n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179,
         n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189,
         n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199,
         n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209,
         n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219,
         n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229,
         n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239,
         n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249,
         n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259,
         n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269,
         n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279,
         n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289,
         n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299,
         n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309,
         n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319,
         n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329,
         n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339,
         n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349,
         n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359,
         n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369,
         n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379,
         n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389,
         n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399,
         n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409,
         n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419,
         n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429,
         n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439,
         n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449,
         n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459,
         n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469,
         n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479,
         n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489,
         n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499,
         n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509,
         n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519,
         n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529,
         n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539,
         n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549,
         n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559,
         n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569,
         n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579,
         n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589,
         n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599,
         n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609,
         n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619,
         n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629,
         n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639,
         n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649,
         n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659,
         n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669,
         n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679,
         n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689,
         n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699,
         n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709,
         n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719,
         n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729,
         n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739,
         n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749,
         n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759,
         n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769,
         n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779,
         n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789,
         n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799,
         n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809,
         n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819,
         n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829,
         n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839,
         n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849,
         n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859,
         n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869,
         n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879,
         n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889,
         n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899,
         n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909,
         n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919,
         n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929,
         n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939,
         n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949,
         n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959,
         n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969,
         n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979,
         n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989,
         n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999,
         n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
         n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
         n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
         n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175,
         n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183,
         n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191,
         n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199,
         n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207,
         n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215,
         n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223,
         n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
         n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239,
         n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247,
         n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255,
         n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263,
         n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271,
         n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279,
         n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287,
         n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295,
         n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303,
         n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311,
         n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319,
         n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327,
         n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335,
         n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343,
         n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351,
         n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359,
         n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367,
         n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375,
         n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383,
         n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391,
         n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399,
         n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407,
         n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415,
         n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423,
         n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431,
         n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439,
         n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447,
         n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455,
         n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463,
         n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471,
         n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479,
         n10480, n10481, n10482, n10483, n10484, n10485, n10486, n10487,
         n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495,
         n10496, n10497, n10498, n10499, n10500, n10501, n10502, n10503,
         n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511,
         n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519,
         n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527,
         n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535,
         n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543,
         n10544, n10545, n10546, n10547, n10548, n10549, n10550, n10551,
         n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559,
         n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567,
         n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575,
         n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583,
         n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591,
         n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599,
         n10600, n10601, n10602, n10603, n10604, n10605, n10606, n10607,
         n10608, n10609, n10610, n10611, n10612, n10613, n10614, n10615,
         n10616, n10617, n10618, n10619, n10620, n10621, n10622, n10623,
         n10624, n10625, n10626, n10627, n10628, n10629, n10630, n10631,
         n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639,
         n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647,
         n10648, n10649, n10650, n10651, n10652, n10653, n10654, n10655,
         n10656, n10657, n10658, n10659, n10660, n10661, n10662, n10663,
         n10664, n10665, n10666, n10667, n10668, n10669, n10670, n10671,
         n10672, n10673, n10674, n10675, n10676, n10677, n10678, n10679,
         n10680, n10681, n10682, n10683, n10684, n10685, n10686, n10687,
         n10688, n10689, n10690, n10691, n10692, n10693, n10694, n10695,
         n10696, n10697, n10698, n10699, n10700, n10701, n10702, n10703,
         n10704, n10705, n10706, n10707, n10708, n10709, n10710, n10711,
         n10712, n10713, n10714, n10715, n10716, n10717, n10718, n10719,
         n10720, n10721, n10722, n10723, n10724, n10725, n10726, n10727,
         n10728, n10729, n10730, n10731, n10732, n10733, n10734, n10735,
         n10736, n10737, n10738, n10739, n10740, n10741, n10742, n10743,
         n10744, n10745, n10746, n10747, n10748, n10749, n10750, n10751,
         n10752, n10753, n10754, n10755, n10756, n10757, n10758, n10759,
         n10760, n10761, n10762, n10763, n10764, n10765, n10766, n10767,
         n10768, n10769, n10770, n10771, n10772, n10773, n10774, n10775,
         n10776, n10777, n10778, n10779, n10780, n10781, n10782, n10783,
         n10784, n10785, n10786, n10787, n10788, n10789, n10790, n10791,
         n10792, n10793, n10794, n10795, n10796, n10797, n10798, n10799,
         n10800, n10801, n10802, n10803, n10804, n10805, n10806, n10807,
         n10808, n10809, n10810, n10811, n10812, n10813, n10814, n10815,
         n10816, n10817, n10818, n10819, n10820, n10821, n10822, n10823,
         n10824, n10825, n10826, n10827, n10828, n10829, n10830, n10831,
         n10832, n10833, n10834, n10835, n10836, n10837, n10838, n10839,
         n10840, n10841, n10842, n10843, n10844, n10845, n10846, n10847,
         n10848, n10849, n10850, n10851, n10852, n10853, n10854, n10855,
         n10856, n10857, n10858, n10859, n10860, n10861, n10862, n10863,
         n10864, n10865, n10866, n10867, n10868, n10869, n10870, n10871,
         n10872, n10873, n10874, n10875, n10876, n10877, n10878, n10879,
         n10880, n10881, n10882, n10883, n10884, n10885, n10886, n10887,
         n10888, n10889, n10890, n10891, n10892, n10893, n10894, n10895,
         n10896, n10897, n10898, n10899, n10900, n10901, n10902, n10903,
         n10904, n10905, n10906, n10907, n10908, n10909, n10910, n10911,
         n10912, n10913, n10914, n10915, n10916, n10917, n10918, n10919,
         n10920, n10921, n10922, n10923, n10924, n10925, n10926, n10927,
         n10928, n10929, n10930, n10931, n10932, n10933, n10934, n10935,
         n10936, n10937, n10938, n10939, n10940, n10941, n10942, n10943,
         n10944, n10945, n10946, n10947, n10948, n10949, n10950, n10951,
         n10952, n10953, n10954, n10955, n10956, n10957, n10958, n10959,
         n10960, n10961, n10962, n10963, n10964, n10965, n10966, n10967,
         n10968, n10969, n10970, n10971, n10972, n10973, n10974, n10975,
         n10976, n10977, n10978, n10979, n10980, n10981, n10982, n10983,
         n10984, n10985, n10986, n10987, n10988, n10989, n10990, n10991,
         n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999,
         n11000, n11001, n11002, n11003, n11004, n11005, n11006, n11007,
         n11008, n11009, n11010, n11011, n11012, n11013, n11014, n11015,
         n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11023,
         n11024, n11025, n11026, n11027, n11028, n11029, n11030, n11031,
         n11032, n11033, n11034, n11035, n11036, n11037, n11038, n11039,
         n11040, n11041, n11042, n11043, n11044, n11045, n11046, n11047,
         n11048, n11049, n11050, n11051, n11052, n11053, n11054, n11055,
         n11056, n11057, n11058, n11059, n11060, n11061, n11062, n11063,
         n11064, n11065, n11066, n11067, n11068, n11069, n11070, n11071,
         n11072, n11073, n11074, n11075, n11076, n11077, n11078, n11079,
         n11080, n11081, n11082, n11083, n11084, n11085, n11086, n11087,
         n11088, n11089, n11090, n11091, n11092, n11093, n11094, n11095,
         n11096, n11097, n11098, n11099, n11100, n11101, n11102, n11103,
         n11104, n11105, n11106, n11107, n11108, n11109, n11110, n11111,
         n11112, n11113, n11114, n11115, n11116, n11117, n11118, n11119,
         n11120, n11121, n11122, n11123, n11124, n11125, n11126, n11127,
         n11128, n11129, n11130, n11131, n11132, n11133, n11134, n11135,
         n11136, n11137, n11138, n11139, n11140, n11141, n11142, n11143,
         n11144, n11145, n11146, n11147, n11148, n11149, n11150, n11151,
         n11152, n11153, n11154, n11155, n11156, n11157, n11158, n11159,
         n11160, n11161, n11162, n11163, n11164, n11165, n11166, n11167,
         n11168, n11169, n11170, n11171, n11172, n11173, n11174, n11175,
         n11176, n11177, n11178, n11179, n11180, n11181, n11182, n11183,
         n11184, n11185, n11186, n11187, n11188, n11189, n11190, n11191,
         n11192, n11193, n11194, n11195, n11196, n11197, n11198, n11199,
         n11200, n11201, n11202, n11203, n11204, n11205, n11206, n11207,
         n11208, n11209, n11210, n11211, n11212, n11213, n11214, n11215,
         n11216, n11217, n11218, n11219, n11220, n11221, n11222, n11223,
         n11224, n11225, n11226, n11227, n11228, n11229, n11230, n11231,
         n11232, n11233, n11234, n11235, n11236, n11237, n11238, n11239,
         n11240, n11241, n11242, n11243, n11244, n11245, n11246, n11247,
         n11248, n11249, n11250, n11251, n11252, n11253, n11254, n11255,
         n11256, n11257, n11258, n11259, n11260, n11261, n11262, n11263,
         n11264, n11265, n11266, n11267, n11268, n11269, n11270, n11271,
         n11272, n11273, n11274, n11275, n11276, n11277, n11278, n11279,
         n11280, n11281, n11282, n11283, n11284, n11285, n11286, n11287,
         n11288, n11289, n11290, n11291, n11292, n11293, n11294, n11295,
         n11296, n11297, n11298, n11299, n11300, n11301, n11302, n11303,
         n11304, n11305, n11306, n11307, n11308, n11309, n11310, n11311,
         n11312, n11313, n11314, n11315, n11316, n11317, n11318, n11319,
         n11320, n11321, n11322, n11323, n11324, n11325, n11326, n11327,
         n11328, n11329, n11330, n11331, n11332, n11333, n11334, n11335,
         n11336, n11337, n11338, n11339, n11340, n11341, n11342, n11343,
         n11344, n11345, n11346, n11347, n11348, n11349, n11350, n11351,
         n11352, n11353, n11354, n11355, n11356, n11357, n11358, n11359,
         n11360, n11361, n11362, n11363, n11364, n11365, n11366, n11367,
         n11368, n11369, n11370, n11371, n11372, n11373, n11374, n11375,
         n11376, n11377, n11378, n11379, n11380, n11381, n11382, n11383,
         n11384, n11385, n11386, n11387, n11388, n11389, n11390, n11391,
         n11392, n11393, n11394, n11395, n11396, n11397, n11398, n11399,
         n11400, n11401, n11402, n11403, n11404, n11405, n11406, n11407,
         n11408, n11409, n11410, n11411, n11412, n11413, n11414, n11415,
         n11416, n11417, n11418, n11419, n11420, n11421, n11422, n11423,
         n11424, n11425, n11426, n11427, n11428, n11429, n11430, n11431,
         n11432, n11433, n11434, n11435, n11436, n11437, n11438, n11439,
         n11440, n11441, n11442, n11443, n11444, n11445, n11446, n11447,
         n11448, n11449, n11450, n11451, n11452, n11453, n11454, n11455,
         n11456, n11457, n11458, n11459, n11460, n11461, n11462, n11463,
         n11464, n11465, n11466, n11467, n11468, n11469, n11470, n11471,
         n11472, n11473, n11474, n11475, n11476, n11477, n11478, n11479,
         n11480, n11481, n11482, n11483, n11484, n11485, n11486, n11487,
         n11488, n11489, n11490, n11491, n11492, n11493, n11494, n11495,
         n11496, n11497, n11498, n11499, n11500, n11501, n11502, n11503,
         n11504, n11505, n11506, n11507, n11508, n11509, n11510, n11511,
         n11512, n11513, n11514, n11515, n11516, n11517, n11518, n11519,
         n11520, n11521, n11522, n11523, n11524, n11525, n11526, n11527,
         n11528, n11529, n11530, n11531, n11532, n11533, n11534, n11535,
         n11536, n11537, n11538, n11539, n11540, n11541, n11542, n11543,
         n11544, n11545, n11546, n11547, n11548, n11549, n11550, n11551,
         n11552, n11553, n11554, n11555, n11556, n11557, n11558, n11559,
         n11560, n11561, n11562, n11563, n11564, n11565, n11566, n11567,
         n11568, n11569, n11570, n11571, n11572, n11573, n11574, n11575,
         n11576, n11577, n11578, n11579, n11580, n11581, n11582, n11583,
         n11584, n11585, n11586, n11587, n11588, n11589, n11590, n11591,
         n11592, n11593, n11594, n11595, n11596, n11597, n11598, n11599,
         n11600, n11601, n11602, n11603, n11604, n11605, n11606, n11607,
         n11608, n11609, n11610, n11611, n11612, n11613, n11614, n11615,
         n11616, n11617, n11618, n11619, n11620, n11621, n11622, n11623,
         n11624, n11625, n11626, n11627, n11628, n11629, n11630, n11631,
         n11632, n11633, n11634, n11635, n11636, n11637, n11638, n11639,
         n11640, n11641, n11642, n11643, n11644, n11645, n11646, n11647,
         n11648, n11649, n11650, n11651, n11652, n11653, n11654, n11655,
         n11656, n11657, n11658, n11659, n11660, n11661, n11662, n11663,
         n11664, n11665, n11666, n11667, n11668, n11669, n11670, n11671,
         n11672, n11673, n11674, n11675, n11676, n11677, n11678, n11679,
         n11680, n11681, n11682, n11683, n11684, n11685, n11686, n11687,
         n11688, n11689, n11690, n11691, n11692, n11693, n11694, n11695,
         n11696, n11697, n11698, n11699, n11700, n11701, n11702, n11703,
         n11704, n11705, n11706, n11707, n11708, n11709, n11710, n11711,
         n11712, n11713, n11714, n11715, n11716, n11717, n11718, n11719,
         n11720, n11721, n11722, n11723, n11724, n11725, n11726, n11727,
         n11728, n11729, n11730, n11731, n11732, n11733, n11734, n11735,
         n11736, n11737, n11738, n11739, n11740, n11741, n11742, n11743,
         n11744, n11745, n11746, n11747, n11748, n11749, n11750, n11751,
         n11752, n11753, n11754, n11755, n11756, n11757, n11758, n11759,
         n11760, n11761, n11762, n11763, n11764, n11765, n11766, n11767,
         n11768, n11769, n11770, n11771, n11772, n11773, n11774, n11775,
         n11776, n11777, n11778, n11779, n11780, n11781, n11782, n11783,
         n11784, n11785, n11786, n11787, n11788, n11789, n11790, n11791,
         n11792, n11793, n11794, n11795, n11796, n11797, n11798, n11799,
         n11800, n11801, n11802, n11803, n11804, n11805, n11806, n11807,
         n11808, n11809, n11810, n11811, n11812, n11813, n11814, n11815,
         n11816, n11817, n11818, n11819, n11820, n11821, n11822, n11823,
         n11824, n11825, n11826, n11827, n11828, n11829, n11830, n11831,
         n11832, n11833, n11834, n11835, n11836, n11837, n11838, n11839,
         n11840, n11841, n11842, n11843, n11844, n11845, n11846, n11847,
         n11848, n11849, n11850, n11851, n11852, n11853, n11854, n11855,
         n11856, n11857, n11858, n11859, n11860, n11861, n11862, n11863,
         n11864, n11865, n11866, n11867, n11868, n11869, n11870, n11871,
         n11872, n11873, n11874, n11875, n11876, n11877, n11878, n11879,
         n11880, n11881, n11882, n11883, n11884, n11885, n11886, n11887,
         n11888, n11889, n11890, n11891, n11892, n11893, n11894, n11895,
         n11896, n11897, n11898, n11899, n11900, n11901, n11902, n11903,
         n11904, n11905, n11906, n11907, n11908, n11909, n11910, n11911,
         n11912, n11913, n11914, n11915, n11916, n11917, n11918, n11919,
         n11920, n11921, n11922, n11923, n11924, n11925, n11926, n11927,
         n11928, n11929, n11930, n11931, n11932, n11933, n11934, n11935,
         n11936, n11937, n11938, n11939, n11940, n11941, n11942, n11943,
         n11944, n11945, n11946, n11947, n11948, n11949, n11950, n11951,
         n11952, n11953, n11954, n11955, n11956, n11957, n11958, n11959,
         n11960, n11961, n11962, n11963, n11964, n11965, n11966, n11967,
         n11968, n11969, n11970, n11971, n11972, n11973, n11974, n11975,
         n11976, n11977, n11978, n11979, n11980, n11981, n11982, n11983,
         n11984, n11985, n11986, n11987, n11988, n11989, n11990, n11991,
         n11992, n11993, n11994, n11995, n11996, n11997, n11998, n11999,
         n12000, n12001, n12002, n12003, n12004, n12005, n12006, n12007,
         n12008, n12009, n12010, n12011, n12012, n12013, n12014, n12015,
         n12016, n12017, n12018, n12019, n12020, n12021, n12022, n12023,
         n12024, n12025, n12026, n12027, n12028, n12029, n12030, n12031,
         n12032, n12033, n12034, n12035, n12036, n12037, n12038, n12039,
         n12040, n12041, n12042, n12043, n12044, n12045, n12046, n12047,
         n12048, n12049, n12050, n12051, n12052, n12053, n12054, n12055,
         n12056, n12057, n12058, n12059, n12060, n12061, n12062, n12063,
         n12064, n12065, n12066, n12067, n12068, n12069, n12070, n12071,
         n12072, n12073, n12074, n12075, n12076, n12077, n12078, n12079,
         n12080, n12081, n12082, n12083, n12084, n12085, n12086, n12087,
         n12088, n12089, n12090, n12091, n12092, n12093, n12094, n12095,
         n12096, n12097, n12098, n12099, n12100, n12101, n12102, n12103,
         n12104, n12105, n12106, n12107, n12108, n12109, n12110, n12111,
         n12112, n12113, n12114, n12115, n12116, n12117, n12118, n12119,
         n12120, n12121, n12122, n12123, n12124, n12125, n12126, n12127,
         n12128, n12129, n12130, n12131, n12132, n12133, n12134, n12135,
         n12136, n12137, n12138, n12139, n12140, n12141, n12142, n12143,
         n12144, n12145, n12146, n12147, n12148, n12149, n12150, n12151,
         n12152, n12153, n12154, n12155, n12156, n12157, n12158, n12159,
         n12160, n12161, n12162, n12163, n12164, n12165, n12166, n12167,
         n12168, n12169, n12170, n12171, n12172, n12173, n12174, n12175,
         n12176, n12177, n12178, n12179, n12180, n12181, n12182, n12183,
         n12184, n12185, n12186, n12187, n12188, n12189, n12190, n12191,
         n12192, n12193, n12194, n12195, n12196, n12197, n12198, n12199,
         n12200, n12201, n12202, n12203, n12204, n12205, n12206, n12207,
         n12208, n12209, n12210, n12211, n12212, n12213, n12214, n12215,
         n12216, n12217, n12218, n12219, n12220, n12221, n12222, n12223,
         n12224, n12225, n12226, n12227, n12228, n12229, n12230, n12231,
         n12232, n12233, n12234, n12235, n12236, n12237, n12238, n12239,
         n12240, n12241, n12242, n12243, n12244, n12245, n12246, n12247,
         n12248, n12249, n12250, n12251, n12252, n12253, n12254, n12255,
         n12256, n12257, n12258, n12259, n12260, n12261, n12262, n12263,
         n12264, n12265, n12266, n12267, n12268, n12269, n12270, n12271,
         n12272, n12273, n12274, n12275, n12276, n12277, n12278, n12279,
         n12280, n12281, n12282, n12283, n12284, n12285, n12286, n12287,
         n12288, n12289, n12290, n12291, n12292, n12293, n12294, n12295,
         n12296, n12297, n12298, n12299, n12300, n12301, n12302, n12303,
         n12304, n12305, n12306, n12307, n12308, n12309, n12310, n12311,
         n12312, n12313, n12314, n12315, n12316, n12317, n12318, n12319,
         n12320, n12321, n12322, n12323, n12324, n12325, n12326, n12327,
         n12328, n12329, n12330, n12331, n12332, n12333, n12334, n12335,
         n12336, n12337, n12338, n12339, n12340, n12341, n12342, n12343,
         n12344, n12345, n12346, n12347, n12348, n12349, n12350, n12351,
         n12352, n12353, n12354, n12355, n12356, n12357, n12358, n12359,
         n12360, n12361, n12362, n12363, n12364, n12365, n12366, n12367,
         n12368, n12369, n12370, n12371, n12372, n12373, n12374, n12375,
         n12376, n12377, n12378, n12379, n12380, n12381, n12382, n12383,
         n12384, n12385, n12386, n12387, n12388, n12389, n12390, n12391,
         n12392, n12393, n12394, n12395, n12396, n12397, n12398, n12399,
         n12400, n12401, n12402, n12403, n12404, n12405, n12406, n12407,
         n12408, n12409, n12410, n12411, n12412, n12413, n12414, n12415,
         n12416, n12417, n12418, n12419, n12420, n12421, n12422, n12423,
         n12424, n12425, n12426, n12427, n12428, n12429, n12430, n12431,
         n12432, n12433, n12434, n12435, n12436, n12437, n12438, n12439,
         n12440, n12441, n12442, n12443, n12444, n12445, n12446, n12447,
         n12448, n12449, n12450, n12451, n12452, n12453, n12454, n12455,
         n12456, n12457, n12458, n12459, n12460, n12461, n12462, n12463,
         n12464, n12465, n12466, n12467, n12468, n12469, n12470, n12471,
         n12472, n12473, n12474, n12475, n12476, n12477, n12478, n12479,
         n12480, n12481, n12482, n12483, n12484, n12485, n12486, n12487,
         n12488, n12489, n12490, n12491, n12492, n12493, n12494, n12495,
         n12496, n12497, n12498, n12499, n12500, n12501, n12502, n12503,
         n12504, n12505, n12506, n12507, n12508, n12509, n12510, n12511,
         n12512, n12513, n12514, n12515, n12516, n12517, n12518, n12519,
         n12520, n12521, n12522, n12523, n12524, n12525, n12526, n12527,
         n12528, n12529, n12530, n12531, n12532, n12533, n12534, n12535,
         n12536, n12537, n12538, n12539, n12540, n12541, n12542, n12543,
         n12544, n12545, n12546, n12547, n12548, n12549, n12550, n12551,
         n12552, n12553, n12554, n12555, n12556, n12557, n12558, n12559,
         n12560, n12561, n12562, n12563, n12564, n12565, n12566, n12567,
         n12568, n12569, n12570, n12571, n12572, n12573, n12574, n12575,
         n12576, n12577, n12578, n12579, n12580, n12581, n12582, n12583,
         n12584, n12585, n12586, n12587, n12588, n12589, n12590, n12591,
         n12592, n12593, n12594, n12595, n12596, n12597, n12598, n12599,
         n12600, n12601, n12602, n12603, n12604, n12605, n12606, n12607,
         n12608, n12609, n12610, n12611, n12612, n12613, n12614, n12615,
         n12616, n12617, n12618, n12619, n12620, n12621, n12622, n12623,
         n12624, n12625, n12626, n12627, n12628, n12629, n12630, n12631,
         n12632, n12633, n12634, n12635, n12636, n12637, n12638, n12639,
         n12640, n12641, n12642, n12643, n12644, n12645, n12646, n12647,
         n12648, n12649, n12650, n12651, n12652, n12653, n12654, n12655,
         n12656, n12657, n12658, n12659, n12660, n12661, n12662, n12663,
         n12664, n12665, n12666, n12667, n12668, n12669, n12670, n12671,
         n12672, n12673, n12674, n12675, n12676, n12677, n12678, n12679,
         n12680, n12681, n12682, n12683, n12684, n12685, n12686, n12687,
         n12688, n12689, n12690, n12691, n12692, n12693, n12694, n12695,
         n12696, n12697, n12698, n12699, n12700, n12701, n12702, n12703,
         n12704, n12705, n12706, n12707, n12708, n12709, n12710, n12711,
         n12712, n12713, n12714, n12715, n12716, n12717, n12718, n12719,
         n12720, n12721, n12722, n12723, n12724, n12725, n12726, n12727,
         n12728, n12729, n12730, n12731, n12732, n12733, n12734, n12735,
         n12736, n12737, n12738, n12739, n12740, n12741, n12742, n12743,
         n12744, n12745, n12746, n12747, n12748, n12749, n12750, n12751,
         n12752, n12753, n12754, n12755, n12756, n12757, n12758, n12759,
         n12760, n12761, n12762, n12763, n12764, n12765, n12766, n12767,
         n12768, n12769, n12770, n12771, n12772, n12773, n12774, n12775,
         n12776, n12777, n12778, n12779, n12780, n12781, n12782, n12783,
         n12784, n12785, n12786, n12787, n12788, n12789, n12790, n12791,
         n12792, n12793, n12794, n12795, n12796, n12797, n12798, n12799,
         n12800, n12801, n12802, n12803, n12804, n12805, n12806, n12807,
         n12808, n12809, n12810, n12811, n12812, n12813, n12814, n12815,
         n12816, n12817, n12818, n12819, n12820, n12821, n12822, n12823,
         n12824, n12825, n12826, n12827, n12828, n12829, n12830, n12831,
         n12832, n12833, n12834, n12835, n12836, n12837, n12838, n12839,
         n12840, n12841, n12842, n12843, n12844, n12845, n12846, n12847,
         n12848, n12849, n12850, n12851, n12852, n12853, n12854, n12855,
         n12856, n12857, n12858, n12859, n12860, n12861, n12862, n12863,
         n12864, n12865, n12866, n12867, n12868, n12869, n12870, n12871,
         n12872, n12873, n12874, n12875, n12876, n12877, n12878, n12879,
         n12880, n12881, n12882, n12883, n12884, n12885, n12886, n12887,
         n12888, n12889, n12890, n12891, n12892, n12893, n12894, n12895,
         n12896, n12897, n12898, n12899, n12900, n12901, n12902, n12903,
         n12904, n12905, n12906, n12907, n12908, n12909, n12910, n12911,
         n12912, n12913, n12914, n12915, n12916, n12917, n12918, n12919,
         n12920, n12921, n12922, n12923, n12924, n12925, n12926, n12927,
         n12928, n12929, n12930, n12931, n12932, n12933, n12934, n12935,
         n12936, n12937, n12938, n12939, n12940, n12941, n12942, n12943,
         n12944, n12945, n12946, n12947, n12948, n12949, n12950, n12951,
         n12952, n12953, n12954, n12955, n12956, n12957, n12958, n12959,
         n12960, n12961, n12962, n12963, n12964, n12965, n12966, n12967,
         n12968, n12969, n12970, n12971, n12972, n12973, n12974, n12975,
         n12976, n12977, n12978, n12979, n12980, n12981, n12982, n12983,
         n12984, n12985, n12986, n12987, n12988, n12989, n12990, n12991,
         n12992, n12993, n12994, n12995, n12996, n12997, n12998, n12999,
         n13000, n13001, n13002, n13003, n13004, n13005, n13006, n13007,
         n13008, n13009, n13010, n13011, n13012, n13013, n13014, n13015,
         n13016, n13017, n13018, n13019, n13020, n13021, n13022, n13023,
         n13024, n13025, n13026, n13027, n13028, n13029, n13030, n13031,
         n13032, n13033, n13034, n13035, n13036, n13037, n13038, n13039,
         n13040, n13041, n13042, n13043, n13044, n13045, n13046, n13047,
         n13048, n13049, n13050, n13051, n13052, n13053, n13054, n13055,
         n13056, n13057, n13058, n13059, n13060, n13061, n13062, n13063,
         n13064, n13065, n13066, n13067, n13068, n13069, n13070, n13071,
         n13072, n13073, n13074, n13075, n13076, n13077, n13078, n13079,
         n13080, n13081, n13082, n13083, n13084, n13085, n13086, n13087,
         n13088, n13089, n13090, n13091, n13092, n13093, n13094, n13095,
         n13096, n13097, n13098, n13099, n13100, n13101, n13102, n13103,
         n13104, n13105, n13106, n13107, n13108, n13109, n13110, n13111,
         n13112, n13113, n13114, n13115, n13116, n13117, n13118, n13119,
         n13120, n13121, n13122, n13123, n13124, n13125, n13126, n13127,
         n13128, n13129, n13130, n13131, n13132, n13133, n13134, n13135,
         n13136, n13137, n13138, n13139, n13140, n13141, n13142, n13143,
         n13144, n13145, n13146, n13147, n13148, n13149, n13150, n13151,
         n13152, n13153, n13154, n13155, n13156, n13157, n13158, n13159,
         n13160, n13161, n13162, n13163, n13164, n13165, n13166, n13167,
         n13168, n13169, n13170, n13171, n13172, n13173, n13174, n13175,
         n13176, n13177, n13178, n13179, n13180, n13181, n13182, n13183,
         n13184, n13185, n13186, n13187, n13188, n13189, n13190, n13191,
         n13192, n13193, n13194, n13195, n13196, n13197, n13198, n13199,
         n13200, n13201, n13202, n13203, n13204, n13205, n13206, n13207,
         n13208, n13209, n13210, n13211, n13212, n13213, n13214, n13215,
         n13216, n13217, n13218, n13219, n13220, n13221, n13222, n13223,
         n13224, n13225, n13226, n13227, n13228, n13229, n13230, n13231,
         n13232, n13233, n13234, n13235, n13236, n13237, n13238, n13239,
         n13240, n13241, n13242, n13243, n13244, n13245, n13246, n13247,
         n13248, n13249, n13250, n13251, n13252, n13253, n13254, n13255,
         n13256, n13257, n13258, n13259, n13260, n13261, n13262, n13263,
         n13264, n13265, n13266, n13267, n13268, n13269, n13270, n13271,
         n13272, n13273, n13274, n13275, n13276, n13277, n13278, n13279,
         n13280, n13281, n13282, n13283, n13284, n13285, n13286, n13287,
         n13288, n13289, n13290, n13291, n13292, n13293, n13294, n13295,
         n13296, n13297, n13298, n13299, n13300, n13301, n13302, n13303,
         n13304, n13305, n13306, n13307, n13308, n13309, n13310, n13311,
         n13312, n13313, n13314, n13315, n13316, n13317, n13318, n13319,
         n13320, n13321, n13322, n13323, n13324, n13325, n13326, n13327,
         n13328, n13329, n13330, n13331, n13332, n13333, n13334, n13335,
         n13336, n13337, n13338, n13339, n13340, n13341, n13342, n13343,
         n13344, n13345, n13346, n13347, n13348, n13349, n13350, n13351,
         n13352, n13353, n13354, n13355, n13356, n13357, n13358, n13359,
         n13360, n13361, n13362, n13363, n13364, n13365, n13366, n13367,
         n13368, n13369, n13370, n13371, n13372, n13373, n13374, n13375,
         n13376, n13377, n13378, n13379, n13380, n13381, n13382, n13383,
         n13384, n13385, n13386, n13387, n13388, n13389, n13390, n13391,
         n13392, n13393, n13394, n13395, n13396, n13397, n13398, n13399,
         n13400, n13401, n13402, n13403, n13404, n13405, n13406, n13407,
         n13408, n13409, n13410, n13411, n13412, n13413, n13414, n13415,
         n13416, n13417, n13418, n13419, n13420, n13421, n13422, n13423,
         n13424, n13425, n13426, n13427, n13428, n13429, n13430, n13431,
         n13432, n13433, n13434, n13435, n13436, n13437, n13438, n13439,
         n13440, n13441, n13442, n13443, n13444, n13445, n13446, n13447,
         n13448, n13449, n13450, n13451, n13452, n13453, n13454, n13455,
         n13456, n13457, n13458, n13459, n13460, n13461, n13462, n13463,
         n13464, n13465, n13466, n13467, n13468, n13469, n13470, n13471,
         n13472, n13473, n13474, n13475, n13476, n13477, n13478, n13479,
         n13480, n13481, n13482, n13483, n13484, n13485, n13486, n13487,
         n13488, n13489, n13490, n13491, n13492, n13493, n13494, n13495,
         n13496, n13497, n13498, n13499, n13500, n13501, n13502, n13503,
         n13504, n13505, n13506, n13507, n13508, n13509, n13510, n13511,
         n13512, n13513, n13514, n13515, n13516, n13517, n13518, n13519,
         n13520, n13521, n13522, n13523, n13524, n13525, n13526, n13527,
         n13528, n13529, n13530, n13531, n13532, n13533, n13534, n13535,
         n13536, n13537, n13538, n13539, n13540, n13541, n13542, n13543,
         n13544, n13545, n13546, n13547, n13548, n13549, n13550, n13551,
         n13552, n13553, n13554, n13555, n13556, n13557, n13558, n13559,
         n13560, n13561, n13562, n13563, n13564, n13565, n13566, n13567,
         n13568, n13569, n13570, n13571, n13572, n13573, n13574, n13575,
         n13576, n13577, n13578, n13579, n13580, n13581, n13582, n13583,
         n13584, n13585, n13586, n13587, n13588, n13589, n13590, n13591,
         n13592, n13593, n13594, n13595, n13596, n13597, n13598, n13599,
         n13600, n13601, n13602, n13603, n13604, n13605, n13606, n13607,
         n13608, n13609, n13610, n13611, n13612, n13613, n13614, n13615,
         n13616, n13617, n13618, n13619, n13620, n13621, n13622, n13623,
         n13624, n13625, n13626, n13627, n13628, n13629, n13630, n13631,
         n13632, n13633, n13634, n13635, n13636, n13637, n13638, n13639,
         n13640, n13641, n13642, n13643, n13644, n13645, n13646, n13647,
         n13648, n13649, n13650, n13651, n13652, n13653, n13654, n13655,
         n13656, n13657, n13658, n13659, n13660, n13661, n13662, n13663,
         n13664, n13665, n13666, n13667, n13668, n13669, n13670, n13671,
         n13672, n13673, n13674, n13675, n13676, n13677, n13678, n13679,
         n13680, n13681, n13682, n13683, n13684, n13685, n13686, n13687,
         n13688, n13689, n13690, n13691, n13692, n13693, n13694, n13695,
         n13696, n13697, n13698, n13699, n13700, n13701, n13702, n13703,
         n13704, n13705, n13706, n13707, n13708, n13709, n13710, n13711,
         n13712, n13713, n13714, n13715, n13716, n13717, n13718, n13719,
         n13720, n13721, n13722, n13723, n13724, n13725, n13726, n13727,
         n13728, n13729, n13730, n13731, n13732, n13733, n13734, n13735,
         n13736, n13737, n13738, n13739, n13740, n13741, n13742, n13743,
         n13744, n13745, n13746, n13747, n13748, n13749, n13750, n13751,
         n13752, n13753, n13754, n13755, n13756, n13757, n13758, n13759,
         n13760, n13761, n13762, n13763, n13764, n13765, n13766, n13767,
         n13768, n13769, n13770, n13771, n13772, n13773, n13774, n13775,
         n13776, n13777, n13778, n13779, n13780, n13781, n13782, n13783,
         n13784, n13785, n13786, n13787, n13788, n13789, n13790, n13791,
         n13792, n13793, n13794, n13795, n13796, n13797, n13798, n13799,
         n13800, n13801, n13802, n13803, n13804, n13805, n13806, n13807,
         n13808, n13809, n13810, n13811, n13812, n13813, n13814, n13815,
         n13816, n13817, n13818, n13819, n13820, n13821, n13822, n13823,
         n13824, n13825, n13826, n13827, n13828, n13829, n13830, n13831,
         n13832, n13833, n13834, n13835, n13836, n13837, n13838, n13839,
         n13840, n13841, n13842, n13843, n13844, n13845, n13846, n13847,
         n13848, n13849, n13850, n13851, n13852, n13853, n13854, n13855,
         n13856, n13857, n13858, n13859, n13860, n13861, n13862, n13863,
         n13864, n13865, n13866, n13867, n13868, n13869, n13870, n13871,
         n13872, n13873, n13874, n13875, n13876, n13877, n13878, n13879,
         n13880, n13881, n13882, n13883, n13884, n13885, n13886, n13887,
         n13888, n13889, n13890, n13891, n13892, n13893, n13894, n13895,
         n13896, n13897, n13898, n13899, n13900, n13901, n13902, n13903,
         n13904, n13905, n13906, n13907, n13908, n13909, n13910, n13911,
         n13912, n13913, n13914, n13915, n13916, n13917, n13918, n13919,
         n13920, n13921, n13922, n13923, n13924, n13925, n13926, n13927,
         n13928, n13929, n13930, n13931, n13932, n13933, n13934, n13935,
         n13936, n13937, n13938, n13939, n13940, n13941, n13942, n13943,
         n13944, n13945, n13946, n13947, n13948, n13949, n13950, n13951,
         n13952, n13953, n13954, n13955, n13956, n13957, n13958, n13959,
         n13960, n13961, n13962, n13963, n13964, n13965, n13966, n13967,
         n13968, n13969, n13970, n13971, n13972, n13973, n13974, n13975,
         n13976, n13977, n13978, n13979, n13980, n13981, n13982, n13983,
         n13984, n13985, n13986, n13987, n13988, n13989, n13990, n13991,
         n13992, n13993, n13994, n13995, n13996, n13997, n13998, n13999,
         n14000, n14001, n14002, n14003, n14004, n14005, n14006, n14007,
         n14008, n14009, n14010, n14011, n14012, n14013, n14014, n14015,
         n14016, n14017, n14018, n14019, n14020, n14021, n14022, n14023,
         n14024, n14025, n14026, n14027, n14028, n14029, n14030, n14031,
         n14032, n14033, n14034, n14035, n14036, n14037, n14038, n14039,
         n14040, n14041, n14042, n14043, n14044, n14045, n14046, n14047,
         n14048, n14049, n14050, n14051, n14052, n14053, n14054, n14055,
         n14056, n14057, n14058, n14059, n14060, n14061, n14062, n14063,
         n14064, n14065, n14066, n14067, n14068, n14069, n14070, n14071,
         n14072, n14073, n14074, n14075, n14076, n14077, n14078, n14079,
         n14080, n14081, n14082, n14083, n14084, n14085, n14086, n14087,
         n14088, n14089, n14090, n14091, n14092, n14093, n14094, n14095,
         n14096, n14097, n14098, n14099, n14100, n14101, n14102, n14103,
         n14104, n14105, n14106, n14107, n14108, n14109, n14110, n14111,
         n14112, n14113, n14114, n14115, n14116, n14117, n14118, n14119,
         n14120, n14121, n14122, n14123, n14124, n14125, n14126, n14127,
         n14128, n14129, n14130, n14131, n14132, n14133, n14134, n14135,
         n14136, n14137, n14138, n14139, n14140, n14141, n14142, n14143,
         n14144, n14145, n14146, n14147, n14148, n14149, n14150, n14151,
         n14152, n14153, n14154, n14155, n14156, n14157, n14158, n14159,
         n14160, n14161, n14162, n14163, n14164, n14165, n14166, n14167,
         n14168, n14169, n14170, n14171, n14172, n14173, n14174, n14175,
         n14176, n14177, n14178, n14179, n14180, n14181, n14182, n14183,
         n14184, n14185, n14186, n14187, n14188, n14189, n14190, n14191,
         n14192, n14193, n14194, n14195, n14196, n14197, n14198, n14199,
         n14200, n14201, n14202, n14203, n14204, n14205, n14206, n14207,
         n14208, n14209, n14210, n14211, n14212, n14213, n14214, n14215,
         n14216, n14217, n14218, n14219, n14220, n14221, n14222, n14223,
         n14224, n14225, n14226, n14227, n14228, n14229, n14230, n14231,
         n14232, n14233, n14234, n14235, n14236, n14237, n14238, n14239,
         n14240, n14241, n14242, n14243, n14244, n14245, n14246, n14247,
         n14248, n14249, n14250, n14251, n14252, n14253, n14254, n14255,
         n14256, n14257, n14258, n14259, n14260, n14261, n14262, n14263,
         n14264, n14265, n14266, n14267, n14268, n14269, n14270, n14271,
         n14272, n14273, n14274, n14275, n14276, n14277, n14278, n14279,
         n14280, n14281, n14282, n14283, n14284, n14285, n14286, n14287,
         n14288, n14289, n14290, n14291, n14292, n14293, n14294, n14295,
         n14296, n14297, n14298, n14299, n14300, n14301, n14302, n14303,
         n14304, n14305, n14306, n14307, n14308, n14309, n14310, n14311,
         n14312, n14313, n14314, n14315, n14316, n14317, n14318, n14319,
         n14320, n14321, n14322, n14323, n14324, n14325, n14326, n14327,
         n14328, n14329, n14330, n14331, n14332, n14333, n14334, n14335,
         n14336, n14337, n14338, n14339, n14340, n14341, n14342, n14343,
         n14344, n14345, n14346, n14347, n14348, n14349, n14350, n14351,
         n14352, n14353, n14354, n14355, n14356, n14357, n14358, n14359,
         n14360, n14361, n14362, n14363, n14364, n14365, n14366, n14367,
         n14368, n14369, n14370, n14371, n14372, n14373, n14374, n14375,
         n14376, n14377, n14378, n14379, n14380, n14381, n14382, n14383,
         n14384, n14385, n14386, n14387, n14388, n14389, n14390, n14391,
         n14392, n14393, n14394, n14395, n14396, n14397, n14398, n14399,
         n14400, n14401, n14402, n14403, n14404, n14405, n14406, n14407,
         n14408, n14409, n14410, n14411, n14412, n14413, n14414, n14415,
         n14416, n14417, n14418, n14419, n14420, n14421, n14422, n14423,
         n14424, n14425, n14426, n14427, n14428, n14429, n14430, n14431,
         n14432, n14433, n14434, n14435, n14436, n14437, n14438, n14439,
         n14440, n14441, n14442, n14443, n14444, n14445, n14446, n14447,
         n14448, n14449, n14450, n14451, n14452, n14453, n14454, n14455,
         n14456, n14457, n14458, n14459, n14460, n14461, n14462, n14463,
         n14464, n14465, n14466, n14467, n14468, n14469, n14470, n14471,
         n14472, n14473, n14474, n14475, n14476, n14477, n14478, n14479,
         n14480, n14481, n14482, n14483, n14484, n14485, n14486, n14487,
         n14488, n14489, n14490, n14491, n14492, n14493, n14494, n14495,
         n14496, n14497, n14498, n14499, n14500, n14501, n14502, n14503,
         n14504, n14505, n14506, n14507, n14508, n14509, n14510, n14511,
         n14512, n14513, n14514, n14515, n14516, n14517, n14518, n14519,
         n14520, n14521, n14522, n14523, n14524, n14525, n14526, n14527,
         n14528, n14529, n14530, n14531, n14532, n14533, n14534, n14535,
         n14536, n14537, n14538, n14539, n14540, n14541, n14542, n14543,
         n14544, n14545, n14546, n14547, n14548, n14549, n14550, n14551,
         n14552, n14553, n14554, n14555, n14556, n14557, n14558, n14559,
         n14560, n14561, n14562, n14563, n14564, n14565, n14566, n14567,
         n14568, n14569, n14570, n14571, n14572, n14573, n14574, n14575,
         n14576, n14577, n14578, n14579, n14580, n14581, n14582, n14583,
         n14584, n14585, n14586, n14587, n14588, n14589, n14590, n14591,
         n14592, n14593, n14594, n14595, n14596, n14597, n14598, n14599,
         n14600, n14601, n14602, n14603, n14604, n14605, n14606, n14607,
         n14608, n14609, n14610, n14611, n14612, n14613, n14614, n14615,
         n14616, n14617, n14618, n14619, n14620, n14621, n14622, n14623,
         n14624, n14625, n14626, n14627, n14628, n14629, n14630, n14631,
         n14632, n14633, n14634, n14635, n14636, n14637, n14638, n14639,
         n14640, n14641, n14642, n14643, n14644, n14645, n14646, n14647,
         n14648, n14649, n14650, n14651, n14652, n14653, n14654, n14655,
         n14656, n14657, n14658, n14659, n14660, n14661, n14662, n14663,
         n14664, n14665, n14666, n14667, n14668, n14669, n14670, n14671,
         n14672, n14673, n14674, n14675, n14676, n14677, n14678, n14679,
         n14680, n14681, n14682, n14683, n14684, n14685, n14686, n14687,
         n14688, n14689, n14690, n14691, n14692, n14693, n14694, n14695,
         n14696, n14697, n14698, n14699, n14700, n14701, n14702, n14703,
         n14704, n14705, n14706, n14707, n14708, n14709, n14710, n14711,
         n14712, n14713, n14714, n14715, n14716, n14717, n14718, n14719,
         n14720, n14721, n14722, n14723, n14724, n14725, n14726, n14727,
         n14728, n14729, n14730, n14731, n14732, n14733, n14734, n14735,
         n14736, n14737, n14738, n14739, n14740, n14741, n14742, n14743,
         n14744, n14745, n14746, n14747, n14748, n14749, n14750, n14751,
         n14752, n14753, n14754, n14755, n14756, n14757, n14758, n14759,
         n14760, n14761, n14762, n14763, n14764, n14765, n14766, n14767,
         n14768, n14769, n14770, n14771, n14772, n14773, n14774, n14775,
         n14776, n14777, n14778, n14779, n14780, n14781, n14782, n14783,
         n14784, n14785, n14786, n14787, n14788, n14789, n14790, n14791,
         n14792, n14793, n14794, n14795, n14796, n14797, n14798, n14799,
         n14800, n14801, n14802, n14803, n14804, n14805, n14806, n14807,
         n14808, n14809, n14810, n14811, n14812, n14813, n14814, n14815,
         n14816, n14817, n14818, n14819, n14820, n14821, n14822, n14823,
         n14824, n14825, n14826, n14827, n14828, n14829, n14830, n14831,
         n14832, n14833, n14834, n14835, n14836, n14837, n14838, n14839,
         n14840, n14841, n14842, n14843, n14844, n14845, n14846, n14847,
         n14848, n14849, n14850, n14851, n14852, n14853, n14854, n14855,
         n14856, n14857, n14858, n14859, n14860, n14861, n14862, n14863,
         n14864, n14865, n14866, n14867, n14868, n14869, n14870, n14871,
         n14872, n14873, n14874, n14875, n14876, n14877, n14878, n14879,
         n14880, n14881, n14882, n14883, n14884, n14885, n14886, n14887,
         n14888, n14889, n14890, n14891, n14892, n14893, n14894, n14895,
         n14896, n14897, n14898, n14899, n14900, n14901, n14902, n14903,
         n14904, n14905, n14906, n14907, n14908, n14909, n14910, n14911,
         n14912, n14913, n14914, n14915, n14916, n14917, n14918, n14919,
         n14920, n14921, n14922, n14923, n14924, n14925, n14926, n14927,
         n14928, n14929, n14930, n14931, n14932, n14933, n14934, n14935,
         n14936, n14937, n14938, n14939, n14940, n14941, n14942, n14943,
         n14944, n14945, n14946, n14947, n14948, n14949, n14950, n14951,
         n14952, n14953, n14954, n14955, n14956, n14957, n14958, n14959,
         n14960, n14961, n14962, n14963, n14964, n14965, n14966, n14967,
         n14968, n14969, n14970, n14971, n14972, n14973, n14974, n14975,
         n14976, n14977, n14978, n14979, n14980, n14981, n14982, n14983,
         n14984, n14985, n14986, n14987, n14988, n14989, n14990, n14991,
         n14992, n14993, n14994, n14995, n14996, n14997, n14998, n14999,
         n15000, n15001, n15002, n15003, n15004, n15005, n15006, n15007,
         n15008, n15009, n15010, n15011, n15012, n15013, n15014, n15015,
         n15016, n15017, n15018, n15019, n15020, n15021, n15022, n15023,
         n15024, n15025, n15026, n15027, n15028, n15029, n15030, n15031,
         n15032, n15033, n15034, n15035, n15036, n15037, n15038, n15039,
         n15040, n15041, n15042, n15043, n15044, n15045, n15046, n15047,
         n15048, n15049, n15050, n15051, n15052, n15053, n15054, n15055,
         n15056, n15057, n15058, n15059, n15060, n15061, n15062, n15063,
         n15064, n15065, n15066, n15067, n15068, n15069, n15070, n15071,
         n15072, n15073, n15074, n15075, n15076, n15077, n15078, n15079,
         n15080, n15081, n15082, n15083, n15084, n15085, n15086, n15087,
         n15088, n15089, n15090, n15091, n15092, n15093, n15094, n15095,
         n15096, n15097, n15098, n15099, n15100, n15101, n15102, n15103,
         n15104, n15105, n15106, n15107, n15108, n15109, n15110, n15111,
         n15112, n15113, n15114, n15115, n15116, n15117, n15118, n15119,
         n15120, n15121, n15122, n15123, n15124, n15125, n15126, n15127,
         n15128, n15129, n15130, n15131, n15132, n15133, n15134, n15135,
         n15136, n15137, n15138, n15139, n15140, n15141, n15142, n15143,
         n15144, n15145, n15146, n15147, n15148, n15149, n15150, n15151,
         n15152, n15153, n15154, n15155, n15156, n15157, n15158, n15159,
         n15160, n15161, n15162, n15163, n15164, n15165, n15166, n15167,
         n15168, n15169, n15170, n15171, n15172, n15173, n15174, n15175,
         n15176, n15177, n15178, n15179, n15180, n15181, n15182, n15183,
         n15184, n15185, n15186, n15187, n15188, n15189, n15190, n15191,
         n15192, n15193, n15194, n15195, n15196, n15197, n15198, n15199,
         n15200, n15201, n15202, n15203, n15204, n15205, n15206, n15207,
         n15208, n15209, n15210, n15211, n15212, n15213, n15214, n15215,
         n15216, n15217, n15218, n15219, n15220, n15221, n15222, n15223,
         n15224, n15225, n15226, n15227, n15228, n15229, n15230, n15231,
         n15232, n15233, n15234, n15235, n15236, n15237, n15238, n15239,
         n15240, n15241, n15242, n15243, n15244, n15245, n15246, n15247,
         n15248, n15249, n15250, n15251, n15252, n15253, n15254, n15255,
         n15256, n15257, n15258, n15259, n15260, n15261, n15262, n15263,
         n15264, n15265, n15266, n15267, n15268, n15269, n15270, n15271,
         n15272, n15273, n15274, n15275, n15276, n15277, n15278, n15279,
         n15280, n15281, n15282, n15283, n15284, n15285, n15286, n15287,
         n15288, n15289, n15290, n15291, n15292, n15293, n15294, n15295,
         n15296, n15297, n15298, n15299, n15300, n15301, n15302, n15303,
         n15304, n15305, n15306, n15307, n15308, n15309, n15310, n15311,
         n15312, n15313, n15314, n15315, n15316, n15317, n15318, n15319,
         n15320, n15321, n15322, n15323, n15324, n15325, n15326, n15327,
         n15328, n15329, n15330, n15331, n15332, n15333, n15334, n15335,
         n15336, n15337, n15338, n15339, n15340, n15341, n15342, n15343,
         n15344, n15345, n15346, n15347, n15348, n15349, n15350, n15351,
         n15352, n15353, n15354, n15355, n15356, n15357, n15358, n15359,
         n15360, n15361, n15362, n15363, n15364, n15365, n15366, n15367,
         n15368, n15369, n15370, n15371, n15372, n15373, n15374, n15375,
         n15376, n15377, n15378, n15379, n15380, n15381, n15382, n15383,
         n15384, n15385, n15386, n15387, n15388, n15389, n15390, n15391,
         n15392, n15393, n15394, n15395, n15396, n15397, n15398, n15399,
         n15400, n15401, n15402, n15403, n15404, n15405, n15406, n15407,
         n15408, n15409, n15410, n15411, n15412, n15413, n15414, n15415,
         n15416, n15417, n15418, n15419, n15420, n15421, n15422, n15423,
         n15424, n15425, n15426, n15427, n15428, n15429, n15430, n15431,
         n15432, n15433, n15434, n15435, n15436, n15437, n15438, n15439,
         n15440, n15441, n15442, n15443, n15444, n15445, n15446, n15447,
         n15448, n15449, n15450, n15451, n15452, n15453, n15454, n15455,
         n15456, n15457, n15458, n15459, n15460, n15461, n15462, n15463,
         n15464, n15465, n15466, n15467, n15468, n15469, n15470, n15471,
         n15472, n15473, n15474, n15475, n15476, n15477, n15478, n15479,
         n15480, n15481, n15482, n15483, n15484, n15485, n15486, n15487,
         n15488, n15489, n15490, n15491, n15492, n15493, n15494, n15495,
         n15496, n15497, n15498, n15499, n15500, n15501, n15502, n15503,
         n15504, n15505, n15506, n15507, n15508, n15509, n15510, n15511,
         n15512, n15513, n15514, n15515, n15516, n15517, n15518, n15519,
         n15520, n15521, n15522, n15523, n15524, n15525, n15526, n15527,
         n15528, n15529, n15530, n15531, n15532, n15533, n15534, n15535,
         n15536, n15537, n15538, n15539, n15540, n15541, n15542, n15543,
         n15544, n15545, n15546, n15547, n15548, n15549, n15550, n15551,
         n15552, n15553, n15554, n15555, n15556, n15557, n15558, n15559,
         n15560, n15561, n15562, n15563, n15564, n15565, n15566, n15567,
         n15568, n15569, n15570, n15571, n15572, n15573, n15574, n15575,
         n15576, n15577, n15578, n15579, n15580, n15581, n15582, n15583,
         n15584, n15585, n15586, n15587, n15588, n15589, n15590, n15591,
         n15592, n15593, n15594, n15595, n15596, n15597, n15598, n15599,
         n15600, n15601, n15602, n15603, n15604, n15605, n15606, n15607,
         n15608, n15609, n15610, n15611, n15612, n15613, n15614, n15615,
         n15616, n15617, n15618, n15619, n15620, n15621, n15622, n15623,
         n15624, n15625, n15626, n15627, n15628, n15629, n15630, n15631,
         n15632, n15633, n15634, n15635, n15636, n15637, n15638, n15639,
         n15640, n15641, n15642, n15643, n15644, n15645, n15646, n15647,
         n15648, n15649, n15650, n15651, n15652, n15653, n15654, n15655,
         n15656, n15657, n15658, n15659, n15660, n15661, n15662, n15663,
         n15664, n15665, n15666, n15667, n15668, n15669, n15670, n15671,
         n15672, n15673, n15674, n15675, n15676, n15677, n15678, n15679,
         n15680, n15681, n15682, n15683, n15684, n15685, n15686, n15687,
         n15688, n15689, n15690, n15691, n15692, n15693, n15694, n15695,
         n15696, n15697, n15698, n15699, n15700, n15701, n15702, n15703,
         n15704, n15705, n15706, n15707, n15708, n15709, n15710, n15711,
         n15712, n15713, n15714, n15715, n15716, n15717, n15718, n15719,
         n15720, n15721, n15722, n15723, n15724, n15725, n15726, n15727,
         n15728, n15729, n15730, n15731, n15732, n15733, n15734, n15735,
         n15736, n15737, n15738, n15739, n15740, n15741, n15742, n15743,
         n15744, n15745, n15746, n15747, n15748, n15749, n15750, n15751,
         n15752, n15753, n15754, n15755, n15756, n15757, n15758, n15759,
         n15760, n15761, n15762, n15763, n15764, n15765, n15766, n15767,
         n15768, n15769, n15770, n15771, n15772, n15773, n15774, n15775,
         n15776, n15777, n15778, n15779, n15780, n15781, n15782, n15783,
         n15784, n15785, n15786, n15787, n15788, n15789, n15790, n15791,
         n15792, n15793, n15794, n15795, n15796, n15797, n15798, n15799,
         n15800, n15801, n15802, n15803, n15804, n15805, n15806, n15807,
         n15808, n15809, n15810, n15811, n15812, n15813, n15814, n15815,
         n15816, n15817, n15818, n15819, n15820, n15821, n15822, n15823,
         n15824, n15825, n15826, n15827, n15828, n15829, n15830, n15831,
         n15832, n15833, n15834, n15835, n15836, n15837, n15838, n15839,
         n15840, n15841, n15842, n15843, n15844, n15845, n15846, n15847,
         n15848, n15849, n15850, n15851, n15852, n15853, n15854, n15855,
         n15856, n15857, n15858, n15859, n15860, n15861, n15862, n15863,
         n15864, n15865, n15866, n15867, n15868, n15869, n15870, n15871,
         n15872, n15873, n15874, n15875, n15876, n15877, n15878, n15879,
         n15880, n15881, n15882, n15883, n15884, n15885, n15886, n15887,
         n15888, n15889, n15890, n15891, n15892, n15893, n15894, n15895,
         n15896, n15897, n15898, n15899, n15900, n15901, n15902, n15903,
         n15904, n15905, n15906, n15907, n15908, n15909, n15910, n15911,
         n15912, n15913, n15914, n15915, n15916, n15917, n15918, n15919,
         n15920, n15921, n15922, n15923, n15924, n15925, n15926, n15927,
         n15928, n15929, n15930, n15931, n15932, n15933, n15934, n15935,
         n15936, n15937, n15938, n15939, n15940, n15941, n15942, n15943,
         n15944, n15945, n15946, n15947, n15948, n15949, n15950, n15951,
         n15952, n15953, n15954, n15955, n15956, n15957, n15958, n15959,
         n15960, n15961, n15962, n15963, n15964, n15965, n15966, n15967,
         n15968, n15969, n15970, n15971, n15972, n15973, n15974, n15975,
         n15976, n15977, n15978, n15979, n15980, n15981, n15982, n15983,
         n15984, n15985, n15986, n15987, n15988, n15989, n15990, n15991,
         n15992, n15993, n15994, n15995, n15996, n15997, n15998, n15999,
         n16000, n16001, n16002, n16003, n16004, n16005, n16006, n16007,
         n16008, n16009, n16010, n16011, n16012, n16013, n16014, n16015,
         n16016, n16017, n16018, n16019, n16020, n16021, n16022, n16023,
         n16024, n16025, n16026, n16027, n16028, n16029, n16030, n16031,
         n16032, n16033, n16034, n16035, n16036, n16037, n16038, n16039,
         n16040, n16041, n16042, n16043, n16044, n16045, n16046, n16047,
         n16048, n16049, n16050, n16051, n16052, n16053, n16054, n16055,
         n16056, n16057, n16058, n16059, n16060, n16061, n16062, n16063,
         n16064, n16065, n16066, n16067, n16068, n16069, n16070, n16071,
         n16072, n16073, n16074, n16075, n16076, n16077, n16078, n16079,
         n16080, n16081, n16082, n16083, n16084, n16085, n16086, n16087,
         n16088, n16089, n16090, n16091, n16092, n16093, n16094, n16095,
         n16096, n16097, n16098, n16099, n16100, n16101, n16102, n16103,
         n16104, n16105, n16106, n16107, n16108, n16109, n16110, n16111,
         n16112, n16113, n16114, n16115, n16116, n16117, n16118, n16119,
         n16120, n16121, n16122, n16123, n16124, n16125, n16126, n16127,
         n16128, n16129, n16130, n16131, n16132, n16133, n16134, n16135,
         n16136, n16137, n16138, n16139, n16140, n16141, n16142, n16143,
         n16144, n16145, n16146, n16147, n16148, n16149, n16150, n16151,
         n16152, n16153, n16154, n16155, n16156, n16157, n16158, n16159,
         n16160, n16161, n16162, n16163, n16164, n16165, n16166, n16167,
         n16168, n16169, n16170, n16171, n16172, n16173, n16174, n16175,
         n16176, n16177, n16178, n16179, n16180, n16181, n16182, n16183,
         n16184, n16185, n16186, n16187, n16188, n16189, n16190, n16191,
         n16192, n16193, n16194, n16195, n16196, n16197, n16198, n16199,
         n16200, n16201, n16202, n16203, n16204, n16205, n16206, n16207,
         n16208, n16209, n16210, n16211, n16212, n16213, n16214, n16215,
         n16216, n16217, n16218, n16219, n16220, n16221, n16222, n16223,
         n16224, n16225, n16226, n16227, n16228, n16229, n16230, n16231,
         n16232, n16233, n16234, n16235, n16236, n16237, n16238, n16239,
         n16240, n16241, n16242, n16243, n16244, n16245, n16246, n16247,
         n16248, n16249, n16250, n16251, n16252, n16253, n16254, n16255,
         n16256, n16257, n16258, n16259, n16260, n16261, n16262, n16263,
         n16264, n16265, n16266, n16267, n16268, n16269, n16270, n16271,
         n16272, n16273, n16274, n16275, n16276, n16277, n16278, n16279,
         n16280, n16281, n16282, n16283, n16284, n16285, n16286, n16287,
         n16288, n16289, n16290, n16291, n16292, n16293, n16294, n16295,
         n16296, n16297, n16298, n16299, n16300, n16301, n16302, n16303,
         n16304, n16305, n16306, n16307, n16308, n16309, n16310, n16311,
         n16312, n16313, n16314, n16315, n16316, n16317, n16318, n16319,
         n16320, n16321, n16322, n16323, n16324, n16325, n16326, n16327,
         n16328, n16329, n16330, n16331, n16332, n16333, n16334, n16335,
         n16336, n16337, n16338, n16339, n16340, n16341, n16342, n16343,
         n16344, n16345, n16346, n16347, n16348, n16349, n16350, n16351,
         n16352, n16353, n16354, n16355, n16356, n16357, n16358, n16359,
         n16360, n16361, n16362, n16363, n16364, n16365, n16366, n16367,
         n16368, n16369, n16370, n16371, n16372, n16373, n16374, n16375,
         n16376, n16377, n16378, n16379, n16380, n16381, n16382, n16383,
         n16384, n16385, n16386, n16387, n16388, n16389, n16390, n16391,
         n16392, n16393, n16394, n16395, n16396, n16397, n16398, n16399,
         n16400, n16401, n16402, n16403, n16404, n16405, n16406, n16407,
         n16408, n16409, n16410, n16411, n16412, n16413, n16414, n16415,
         n16416, n16417, n16418, n16419, n16420, n16421, n16422, n16423,
         n16424, n16425, n16426, n16427, n16428, n16429, n16430, n16431,
         n16432, n16433, n16434, n16435, n16436, n16437, n16438, n16439,
         n16440, n16441, n16442, n16443, n16444, n16445, n16446, n16447,
         n16448, n16449, n16450, n16451, n16452, n16453, n16454, n16455,
         n16456, n16457, n16458, n16459, n16460, n16461, n16462, n16463,
         n16464, n16465, n16466, n16467, n16468, n16469, n16470, n16471,
         n16472, n16473, n16474, n16475, n16476, n16477, n16478, n16479,
         n16480, n16481, n16482, n16483, n16484, n16485, n16486, n16487,
         n16488, n16489, n16490, n16491, n16492, n16493, n16494, n16495,
         n16496, n16497, n16498, n16499, n16500, n16501, n16502, n16503,
         n16504, n16505, n16506, n16507, n16508, n16509, n16510, n16511,
         n16512, n16513, n16514, n16515, n16516, n16517, n16518, n16519,
         n16520, n16521, n16522, n16523, n16524, n16525, n16526, n16527,
         n16528, n16529, n16530, n16531, n16532, n16533, n16534, n16535,
         n16536, n16537, n16538, n16539, n16540, n16541, n16542, n16543,
         n16544, n16545, n16546, n16547, n16548, n16549, n16550, n16551,
         n16552, n16553, n16554, n16555, n16556, n16557, n16558, n16559,
         n16560, n16561, n16562, n16563, n16564, n16565, n16566, n16567,
         n16568, n16569, n16570, n16571, n16572, n16573, n16574, n16575,
         n16576, n16577, n16578, n16579, n16580, n16581, n16582, n16583,
         n16584, n16585, n16586, n16587, n16588, n16589, n16590, n16591,
         n16592, n16593, n16594, n16595, n16596, n16597, n16598, n16599,
         n16600, n16601, n16602, n16603, n16604, n16605, n16606, n16607,
         n16608, n16609, n16610, n16611, n16612, n16613, n16614, n16615,
         n16616, n16617, n16618, n16619, n16620, n16621, n16622, n16623,
         n16624, n16625, n16626, n16627, n16628, n16629, n16630, n16631,
         n16632, n16633, n16634, n16635, n16636, n16637, n16638, n16639,
         n16640, n16641, n16642, n16643, n16644, n16645, n16646, n16647,
         n16648, n16649, n16650, n16651, n16652, n16653, n16654, n16655,
         n16656, n16657, n16658, n16659, n16660, n16661, n16662, n16663,
         n16664, n16665, n16666, n16667, n16668, n16669, n16670, n16671,
         n16672, n16673, n16674, n16675, n16676, n16677, n16678, n16679,
         n16680, n16681, n16682, n16683, n16684, n16685, n16686, n16687,
         n16688, n16689, n16690, n16691, n16692, n16693, n16694, n16695,
         n16696, n16697, n16698, n16699, n16700, n16701, n16702, n16703,
         n16704, n16705, n16706, n16707, n16708, n16709, n16710, n16711,
         n16712, n16713, n16714, n16715, n16716, n16717, n16718, n16719,
         n16720, n16721, n16722, n16723, n16724, n16725, n16726, n16727,
         n16728, n16729, n16730, n16731, n16732, n16733, n16734, n16735,
         n16736, n16737, n16738, n16739, n16740, n16741, n16742, n16743,
         n16744, n16745, n16746, n16747, n16748, n16749, n16750, n16751,
         n16752, n16753, n16754, n16755, n16756, n16757, n16758, n16759,
         n16760, n16761, n16762, n16763, n16764, n16765, n16766, n16767,
         n16768, n16769, n16770, n16771, n16772, n16773, n16774, n16775,
         n16776, n16777, n16778, n16779, n16780, n16781, n16782, n16783,
         n16784, n16785, n16786, n16787, n16788, n16789, n16790, n16791,
         n16792, n16793, n16794, n16795, n16796, n16797, n16798, n16799,
         n16800, n16801, n16802, n16803, n16804, n16805, n16806, n16807,
         n16808, n16809, n16810, n16811, n16812, n16813, n16814, n16815,
         n16816, n16817, n16818, n16819, n16820, n16821, n16822, n16823,
         n16824, n16825, n16826, n16827, n16828, n16829, n16830, n16831,
         n16832, n16833, n16834, n16835, n16836, n16837, n16838, n16839,
         n16840, n16841, n16842, n16843, n16844, n16845, n16846, n16847,
         n16848, n16849, n16850, n16851, n16852, n16853, n16854, n16855,
         n16856, n16857, n16858, n16859, n16860, n16861, n16862, n16863,
         n16864, n16865, n16866, n16867, n16868, n16869, n16870, n16871,
         n16872, n16873, n16874, n16875, n16876, n16877, n16878, n16879,
         n16880, n16881, n16882, n16883, n16884, n16885, n16886, n16887,
         n16888, n16889, n16890, n16891, n16892, n16893, n16894, n16895,
         n16896, n16897, n16898, n16899, n16900, n16901, n16902, n16903,
         n16904, n16905, n16906, n16907, n16908, n16909, n16910, n16911,
         n16912, n16913, n16914, n16915, n16916, n16917, n16918, n16919,
         n16920, n16921, n16922, n16923, n16924, n16925, n16926, n16927,
         n16928, n16929, n16930, n16931, n16932, n16933, n16934, n16935,
         n16936, n16937, n16938, n16939, n16940, n16941, n16942, n16943,
         n16944, n16945, n16946, n16947, n16948, n16949, n16950, n16951,
         n16952, n16953, n16954, n16955, n16956, n16957, n16958, n16959,
         n16960, n16961, n16962, n16963, n16964, n16965, n16966, n16967,
         n16968, n16969, n16970, n16971, n16972, n16973, n16974, n16975,
         n16976, n16977, n16978, n16979, n16980, n16981, n16982, n16983,
         n16984, n16985, n16986, n16987, n16988, n16989, n16990, n16991,
         n16992, n16993, n16994, n16995, n16996, n16997, n16998, n16999,
         n17000, n17001, n17002, n17003, n17004, n17005, n17006, n17007,
         n17008, n17009, n17010, n17011, n17012, n17013, n17014, n17015,
         n17016, n17017, n17018, n17019, n17020, n17021, n17022, n17023,
         n17024, n17025, n17026, n17027, n17028, n17029, n17030, n17031,
         n17032, n17033, n17034, n17035, n17036, n17037, n17038, n17039,
         n17040, n17041, n17042, n17043, n17044, n17045, n17046, n17047,
         n17048, n17049, n17050, n17051, n17052, n17053, n17054, n17055,
         n17056, n17057, n17058, n17059, n17060, n17061, n17062, n17063,
         n17064, n17065, n17066, n17067, n17068, n17069, n17070, n17071,
         n17072, n17073, n17074, n17075, n17076, n17077, n17078, n17079,
         n17080, n17081, n17082, n17083, n17084, n17085, n17086, n17087,
         n17088, n17089, n17090, n17091, n17092, n17093, n17094, n17095,
         n17096, n17097, n17098, n17099, n17100, n17101, n17102, n17103,
         n17104, n17105, n17106, n17107, n17108, n17109, n17110, n17111,
         n17112, n17113, n17114, n17115, n17116, n17117, n17118, n17119,
         n17120, n17121, n17122, n17123, n17124, n17125, n17126, n17127,
         n17128, n17129, n17130, n17131, n17132, n17133, n17134, n17135,
         n17136, n17137, n17138, n17139, n17140, n17141, n17142, n17143,
         n17144, n17145, n17146, n17147, n17148, n17149, n17150, n17151,
         n17152, n17153, n17154, n17155, n17156, n17157, n17158, n17159,
         n17160, n17161, n17162, n17163, n17164, n17165, n17166, n17167,
         n17168, n17169, n17170, n17171, n17172, n17173, n17174, n17175,
         n17176, n17177, n17178, n17179, n17180, n17181, n17182, n17183,
         n17184, n17185, n17186, n17187, n17188, n17189, n17190, n17191,
         n17192, n17193, n17194, n17195, n17196, n17197, n17198, n17199,
         n17200, n17201, n17202, n17203, n17204, n17205, n17206, n17207,
         n17208, n17209, n17210, n17211, n17212, n17213, n17214, n17215,
         n17216, n17217, n17218, n17219, n17220, n17221, n17222, n17223,
         n17224, n17225, n17226, n17227, n17228, n17229, n17230, n17231,
         n17232, n17233, n17234, n17235, n17236, n17237, n17238, n17239,
         n17240, n17241, n17242, n17243, n17244, n17245, n17246, n17247,
         n17248, n17249, n17250, n17251, n17252, n17253, n17254, n17255,
         n17256, n17257, n17258, n17259, n17260, n17261, n17262, n17263,
         n17264, n17265, n17266, n17267, n17268, n17269, n17270, n17271,
         n17272, n17273, n17274, n17275, n17276, n17277, n17278, n17279,
         n17280, n17281, n17282, n17283, n17284, n17285, n17286, n17287,
         n17288, n17289, n17290, n17291, n17292, n17293, n17294, n17295,
         n17296, n17297, n17298, n17299, n17300, n17301, n17302, n17303,
         n17304, n17305, n17306, n17307, n17308, n17309, n17310, n17311,
         n17312, n17313, n17314, n17315, n17316, n17317, n17318, n17319,
         n17320, n17321, n17322, n17323, n17324, n17325, n17326, n17327,
         n17328, n17329, n17330, n17331, n17332, n17333, n17334, n17335,
         n17336, n17337, n17338, n17339, n17340, n17341, n17342, n17343,
         n17344, n17345, n17346, n17347, n17348, n17349, n17350, n17351,
         n17352, n17353, n17354, n17355, n17356, n17357, n17358, n17359,
         n17360, n17361, n17362, n17363, n17364, n17365, n17366, n17367,
         n17368, n17369, n17370, n17371, n17372, n17373, n17374, n17375,
         n17376, n17377, n17378, n17379, n17380, n17381, n17382, n17383,
         n17384, n17385, n17386, n17387, n17388, n17389, n17390, n17391,
         n17392, n17393, n17394, n17395, n17396, n17397, n17398, n17399,
         n17400, n17401, n17402, n17403, n17404, n17405, n17406, n17407,
         n17408, n17409, n17410, n17411, n17412, n17413, n17414, n17415,
         n17416, n17417, n17418, n17419, n17420, n17421, n17422, n17423,
         n17424, n17425, n17426, n17427, n17428, n17429, n17430, n17431,
         n17432, n17433, n17434, n17435, n17436, n17437, n17438, n17439,
         n17440, n17441, n17442, n17443, n17444, n17445, n17446, n17447,
         n17448, n17449, n17450, n17451, n17452, n17453, n17454, n17455,
         n17456, n17457, n17458, n17459, n17460, n17461, n17462, n17463,
         n17464, n17465, n17466, n17467, n17468, n17469, n17470, n17471,
         n17472, n17473, n17474, n17475, n17476, n17477, n17478, n17479,
         n17480, n17481, n17482, n17483, n17484, n17485, n17486, n17487,
         n17488, n17489, n17490, n17491, n17492, n17493, n17494, n17495,
         n17496, n17497, n17498, n17499, n17500, n17501, n17502, n17503,
         n17504, n17505, n17506, n17507, n17508, n17509, n17510, n17511,
         n17512, n17513, n17514, n17515, n17516, n17517, n17518, n17519,
         n17520, n17521, n17522, n17523, n17524, n17525, n17526, n17527,
         n17528, n17529, n17530, n17531, n17532, n17533, n17534, n17535,
         n17536, n17537, n17538, n17539, n17540, n17541, n17542, n17543,
         n17544, n17545, n17546, n17547, n17548, n17549, n17550, n17551,
         n17552, n17553, n17554, n17555, n17556, n17557, n17558, n17559,
         n17560, n17561, n17562, n17563, n17564, n17565, n17566, n17567,
         n17568, n17569, n17570, n17571, n17572, n17573, n17574, n17575,
         n17576, n17577, n17578, n17579, n17580, n17581, n17582, n17583,
         n17584, n17585, n17586, n17587, n17588, n17589, n17590, n17591,
         n17592, n17593, n17594, n17595, n17596, n17597, n17598, n17599,
         n17600, n17601, n17602, n17603, n17604, n17605, n17606, n17607,
         n17608, n17609, n17610, n17611, n17612, n17613, n17614, n17615,
         n17616, n17617, n17618, n17619, n17620, n17621, n17622, n17623,
         n17624, n17625, n17626, n17627, n17628, n17629, n17630, n17631,
         n17632, n17633, n17634, n17635, n17636, n17637, n17638, n17639,
         n17640, n17641, n17642, n17643, n17644, n17645, n17646, n17647,
         n17648, n17649, n17650, n17651, n17652, n17653, n17654, n17655,
         n17656, n17657, n17658, n17659, n17660, n17661, n17662, n17663,
         n17664, n17665, n17666, n17667, n17668, n17669, n17670, n17671,
         n17672, n17673, n17674, n17675, n17676, n17677, n17678, n17679,
         n17680, n17681, n17682, n17683, n17684, n17685, n17686, n17687,
         n17688, n17689, n17690, n17691, n17692, n17693, n17694, n17695,
         n17696, n17697, n17698, n17699, n17700, n17701, n17702, n17703,
         n17704, n17705, n17706, n17707, n17708, n17709, n17710, n17711,
         n17712, n17713, n17714, n17715, n17716, n17717, n17718, n17719,
         n17720, n17721, n17722, n17723, n17724, n17725, n17726, n17727,
         n17728, n17729, n17730, n17731, n17732, n17733, n17734, n17735,
         n17736, n17737, n17738, n17739, n17740, n17741, n17742, n17743,
         n17744, n17745, n17746, n17747, n17748, n17749, n17750, n17751,
         n17752, n17753, n17754, n17755, n17756, n17757, n17758, n17759,
         n17760, n17761, n17762, n17763, n17764, n17765, n17766, n17767,
         n17768, n17769, n17770, n17771, n17772, n17773, n17774, n17775,
         n17776, n17777, n17778, n17779, n17780, n17781, n17782, n17783,
         n17784, n17785, n17786, n17787, n17788, n17789, n17790, n17791,
         n17792, n17793, n17794, n17795, n17796, n17797, n17798, n17799,
         n17800, n17801, n17802, n17803, n17804, n17805, n17806, n17807,
         n17808, n17809, n17810, n17811, n17812, n17813, n17814, n17815,
         n17816, n17817, n17818, n17819, n17820, n17821, n17822, n17823,
         n17824, n17825, n17826, n17827, n17828, n17829, n17830, n17831,
         n17832, n17833, n17834, n17835, n17836, n17837, n17838, n17839,
         n17840, n17841, n17842, n17843, n17844, n17845, n17846, n17847,
         n17848, n17849, n17850, n17851, n17852, n17853, n17854, n17855,
         n17856, n17857, n17858, n17859, n17860, n17861, n17862, n17863,
         n17864, n17865, n17866, n17867, n17868, n17869, n17870, n17871,
         n17872, n17873, n17874, n17875, n17876, n17877, n17878, n17879,
         n17880, n17881, n17882, n17883, n17884, n17885, n17886, n17887,
         n17888, n17889, n17890, n17891, n17892, n17893, n17894, n17895,
         n17896, n17897, n17898, n17899, n17900, n17901, n17902, n17903,
         n17904, n17905, n17906, n17907, n17908, n17909, n17910, n17911,
         n17912, n17913, n17914, n17915, n17916, n17917, n17918, n17919,
         n17920, n17921, n17922, n17923, n17924, n17925, n17926, n17927,
         n17928, n17929, n17930, n17931, n17932, n17933, n17934, n17935,
         n17936, n17937, n17938, n17939, n17940, n17941, n17942, n17943,
         n17944, n17945, n17946, n17947, n17948, n17949, n17950, n17951,
         n17952, n17953, n17954, n17955, n17956, n17957, n17958, n17959,
         n17960, n17961, n17962, n17963, n17964, n17965, n17966, n17967,
         n17968, n17969, n17970, n17971, n17972, n17973, n17974, n17975,
         n17976, n17977, n17978, n17979, n17980, n17981, n17982, n17983,
         n17984, n17985, n17986, n17987, n17988, n17989, n17990, n17991,
         n17992, n17993, n17994, n17995, n17996, n17997, n17998, n17999,
         n18000, n18001, n18002, n18003, n18004, n18005, n18006, n18007,
         n18008, n18009, n18010, n18011, n18012, n18013, n18014, n18015,
         n18016, n18017, n18018, n18019, n18020, n18021, n18022, n18023,
         n18024, n18025, n18026, n18027, n18028, n18029, n18030, n18031,
         n18032, n18033, n18034, n18035, n18036, n18037, n18038, n18039,
         n18040, n18041, n18042, n18043, n18044, n18045, n18046, n18047,
         n18048, n18049, n18050, n18051, n18052, n18053, n18054, n18055,
         n18056, n18057, n18058, n18059, n18060, n18061, n18062, n18063,
         n18064, n18065, n18066, n18067, n18068, n18069, n18070, n18071,
         n18072, n18073, n18074, n18075, n18076, n18077, n18078, n18079,
         n18080, n18081, n18082, n18083, n18084, n18085, n18086, n18087,
         n18088, n18089, n18090, n18091, n18092, n18093, n18094, n18095,
         n18096, n18097, n18098, n18099, n18100, n18101, n18102, n18103,
         n18104, n18105, n18106, n18107, n18108, n18109, n18110, n18111,
         n18112, n18113, n18114, n18115, n18116, n18117, n18118, n18119,
         n18120, n18121, n18122, n18123, n18124, n18125, n18126, n18127,
         n18128, n18129, n18130, n18131, n18132, n18133, n18134, n18135,
         n18136, n18137, n18138, n18139, n18140, n18141, n18142, n18143,
         n18144, n18145, n18146, n18147, n18148, n18149, n18150, n18151,
         n18152, n18153, n18154, n18155, n18156, n18157, n18158, n18159,
         n18160, n18161, n18162, n18163, n18164, n18165, n18166, n18167,
         n18168, n18169, n18170, n18171, n18172, n18173, n18174, n18175,
         n18176, n18177, n18178, n18179, n18180, n18181, n18182, n18183,
         n18184, n18185, n18186, n18187, n18188, n18189, n18190, n18191,
         n18192, n18193, n18194, n18195, n18196, n18197, n18198, n18199,
         n18200, n18201, n18202, n18203, n18204, n18205, n18206, n18207,
         n18208, n18209, n18210, n18211, n18212, n18213, n18214, n18215,
         n18216, n18217, n18218, n18219, n18220, n18221, n18222, n18223,
         n18224, n18225, n18226, n18227, n18228, n18229, n18230, n18231,
         n18232, n18233, n18234, n18235, n18236, n18237, n18238, n18239,
         n18240, n18241, n18242, n18243, n18244, n18245, n18246, n18247,
         n18248, n18249, n18250, n18251, n18252, n18253, n18254, n18255,
         n18256, n18257, n18258, n18259, n18260, n18261, n18262, n18263,
         n18264, n18265, n18266, n18267, n18268, n18269, n18270, n18271,
         n18272, n18273, n18274, n18275, n18276, n18277, n18278, n18279,
         n18280, n18281, n18282, n18283, n18284, n18285, n18286, n18287,
         n18288, n18289, n18290, n18291, n18292, n18293, n18294, n18295,
         n18296, n18297, n18298, n18299, n18300, n18301, n18302, n18303,
         n18304, n18305, n18306, n18307, n18308, n18309, n18310, n18311,
         n18312, n18313, n18314, n18315, n18316, n18317, n18318, n18319,
         n18320, n18321, n18322, n18323, n18324, n18325, n18326, n18327,
         n18328, n18329, n18330, n18331, n18332, n18333, n18334, n18335,
         n18336, n18337, n18338, n18339, n18340, n18341, n18342, n18343,
         n18344, n18345, n18346, n18347, n18348, n18349, n18350, n18351,
         n18352, n18353, n18354, n18355, n18356, n18357, n18358, n18359,
         n18360, n18361, n18362, n18363, n18364, n18365, n18366, n18367,
         n18368, n18369, n18370, n18371, n18372, n18373, n18374, n18375,
         n18376, n18377, n18378, n18379, n18380, n18381, n18382, n18383,
         n18384, n18385, n18386, n18387, n18388, n18389, n18390, n18391,
         n18392, n18393, n18394, n18395, n18396, n18397, n18398, n18399,
         n18400, n18401, n18402;
  wire   [219:0] Poly0;
  wire   [219:0] poly0_shifted;
  wire   [346:0] Poly1;
  wire   [346:0] poly1_shifted;
  wire   [69:0] Poly2;
  wire   [69:0] poly2_shifted;
  wire   [83:0] Poly3;
  wire   [83:0] poly3_shifted;
  wire   [60:0] Poly4;
  wire   [60:0] poly4_shifted;
  wire   [124:0] Poly5;
  wire   [124:0] poly5_shifted;
  wire   [55:0] Poly6;
  wire   [55:0] poly6_shifted;
  wire   [410:0] Poly7;
  wire   [410:0] poly7_shifted;
  wire   [95:0] Poly8;
  wire   [95:0] poly8_shifted;
  wire   [115:0] Poly9;
  wire   [115:0] poly9_shifted;
  wire   [42:0] Poly10;
  wire   [42:0] poly10_shifted;
  wire   [85:0] Poly11;
  wire   [85:0] poly11_shifted;
  wire   [126:0] Poly12;
  wire   [126:0] poly12_shifted;
  wire   [527:0] Poly13;
  wire   [527:0] poly13_shifted;
  wire   [300:0] Poly14;
  wire   [300:0] poly14_shifted;
  wire   [59:0] Poly15;
  wire   [59:0] poly15_shifted;
  wire   [15:0] polydata;
  wire   [31:0] scrambler;
  wire   [63:0] dataselector;

  CFD2QX1 \Poly4_reg[60]  ( .D(n8796), .CP(clk), .CD(n18389), .Q(Poly4[60]) );
  CFD2QX1 \Poly4_reg[57]  ( .D(n8799), .CP(clk), .CD(n18256), .Q(Poly4[57]) );
  CFD2QX1 \Poly4_reg[52]  ( .D(n8804), .CP(clk), .CD(n18256), .Q(Poly4[52]) );
  CFD2QX1 \Poly4_reg[59]  ( .D(n8797), .CP(clk), .CD(n18389), .Q(Poly4[59]) );
  CFD2QX1 \Poly4_reg[50]  ( .D(n8806), .CP(clk), .CD(n18389), .Q(Poly4[50]) );
  CFD2QX1 \Poly4_reg[56]  ( .D(n8800), .CP(clk), .CD(n18385), .Q(Poly4[56]) );
  CFD2QX1 \Poly4_reg[54]  ( .D(n8802), .CP(clk), .CD(n18386), .Q(Poly4[54]) );
  CFD2QX1 \dataselector_reg[21]  ( .D(n8774), .CP(clk), .CD(n18402), .Q(
        dataselector[21]) );
  CFD2QX1 \dataselector_reg[63]  ( .D(n8732), .CP(clk), .CD(n18402), .Q(
        dataselector[63]) );
  CFD2QX1 \dataselector_reg[62]  ( .D(n8733), .CP(clk), .CD(n18402), .Q(
        dataselector[62]) );
  CFD2QX1 \dataselector_reg[59]  ( .D(n8736), .CP(clk), .CD(n18402), .Q(
        dataselector[59]) );
  CFD2QX1 \dataselector_reg[58]  ( .D(n8737), .CP(clk), .CD(n18402), .Q(
        dataselector[58]) );
  CFD2QX1 \scrambler_reg[28]  ( .D(n8728), .CP(clk), .CD(n18257), .Q(
        scrambler[28]) );
  CFD2QX1 \scrambler_reg[24]  ( .D(n8724), .CP(clk), .CD(n18257), .Q(
        scrambler[24]) );
  CFD2QX1 \scrambler_reg[22]  ( .D(n8722), .CP(clk), .CD(n18257), .Q(
        scrambler[22]) );
  CFD2QX1 \scrambler_reg[21]  ( .D(n8721), .CP(clk), .CD(n18257), .Q(
        scrambler[21]) );
  CFD2QX1 \scrambler_reg[18]  ( .D(n8718), .CP(clk), .CD(n18257), .Q(
        scrambler[18]) );
  CFD2QX1 \dataselector_reg[14]  ( .D(n8781), .CP(clk), .CD(n18402), .Q(
        dataselector[14]) );
  CFD2QXL \scrambler_reg[26]  ( .D(n8726), .CP(clk), .CD(n18257), .Q(
        scrambler[26]) );
  CFD2QXL \scrambler_reg[9]  ( .D(n8709), .CP(clk), .CD(n18257), .Q(
        scrambler[9]) );
  CFD2QXL \scrambler_reg[17]  ( .D(n8717), .CP(clk), .CD(n18257), .Q(
        scrambler[17]) );
  CFD2QXL \polydata_reg[3]  ( .D(n8687), .CP(clk), .CD(n18257), .Q(polydata[3]) );
  CFD2QXL \polydata_reg[14]  ( .D(n8698), .CP(clk), .CD(n18257), .Q(
        polydata[14]) );
  CFD2QXL \scrambler_reg[12]  ( .D(n8712), .CP(clk), .CD(n18257), .Q(
        scrambler[12]) );
  CFD2QXL \Poly5_reg[24]  ( .D(n11502), .CP(clk), .CD(n18257), .Q(
        poly5_shifted[38]) );
  CFD2QXL \Poly10_reg[1]  ( .D(n11102), .CP(clk), .CD(n18262), .Q(Poly10[1])
         );
  CFD2QXL \Poly1_reg[25]  ( .D(n9332), .CP(clk), .CD(n18361), .Q(Poly1[25]) );
  CFD2QXL \Poly0_reg[206]  ( .D(n9371), .CP(clk), .CD(n18348), .Q(Poly0[206])
         );
  CFD2QXL \Poly5_reg[119]  ( .D(n11407), .CP(clk), .CD(n18259), .Q(Poly5[119])
         );
  CFD2QXL \Poly1_reg[341]  ( .D(n9016), .CP(clk), .CD(n18393), .Q(Poly1[341])
         );
  CFD2QXL \Poly8_reg[90]  ( .D(n11311), .CP(clk), .CD(n18261), .Q(Poly8[90])
         );
  CFD2QXL \Poly6_reg[55]  ( .D(n9638), .CP(clk), .CD(n18342), .Q(Poly6[55]) );
  CFD2QXL \Poly10_reg[35]  ( .D(n11068), .CP(clk), .CD(n18262), .Q(Poly10[35])
         );
  CFD2QXL \Poly5_reg[84]  ( .D(n11442), .CP(clk), .CD(n18257), .Q(Poly5[84])
         );
  CFD2QXL pushin_1d_reg ( .D(n16435), .CP(clk), .CD(n18257), .Q(pushout) );
  CFD2QXL \Poly0_reg[87]  ( .D(n9490), .CP(clk), .CD(n18394), .Q(
        poly0_shifted[105]) );
  CFD2QXL \Poly0_reg[96]  ( .D(n9481), .CP(clk), .CD(n18357), .Q(
        poly0_shifted[114]) );
  CFD2QXL \Poly5_reg[45]  ( .D(n11481), .CP(clk), .CD(n18257), .Q(
        poly5_shifted[59]) );
  CFD2QXL \Poly0_reg[95]  ( .D(n9482), .CP(clk), .CD(n18351), .Q(
        poly0_shifted[113]) );
  CFD2QXL \Poly0_reg[82]  ( .D(n9495), .CP(clk), .CD(n18351), .Q(
        poly0_shifted[100]) );
  CFD2QXL \Poly0_reg[85]  ( .D(n9492), .CP(clk), .CD(n18354), .Q(
        poly0_shifted[103]) );
  CFD2QXL \Poly0_reg[92]  ( .D(n9485), .CP(clk), .CD(n18355), .Q(
        poly0_shifted[110]) );
  CFD2QXL \Poly0_reg[94]  ( .D(n9483), .CP(clk), .CD(n18356), .Q(
        poly0_shifted[112]) );
  CFD2QXL \Poly1_reg[20]  ( .D(n9337), .CP(clk), .CD(n18368), .Q(Poly1[20]) );
  CFD2QXL \dataselector_reg[51]  ( .D(n8744), .CP(clk), .CD(n18257), .Q(
        dataselector[51]) );
  CFD2QXL \polydata_reg[7]  ( .D(n8691), .CP(clk), .CD(n18257), .Q(polydata[7]) );
  CFD2QXL \polydata_reg[9]  ( .D(n8693), .CP(clk), .CD(n18401), .Q(polydata[9]) );
  CFD2QXL \polydata_reg[10]  ( .D(n8694), .CP(clk), .CD(n18257), .Q(
        polydata[10]) );
  CFD2QXL \polydata_reg[8]  ( .D(n8692), .CP(clk), .CD(n18257), .Q(polydata[8]) );
  CFD2QXL \polydata_reg[1]  ( .D(n8685), .CP(clk), .CD(n18257), .Q(polydata[1]) );
  CFD2QXL \polydata_reg[6]  ( .D(n8690), .CP(clk), .CD(n18401), .Q(polydata[6]) );
  CFD2QXL \Poly0_reg[183]  ( .D(n9394), .CP(clk), .CD(n18393), .Q(
        poly0_shifted[201]) );
  CFD2QXL \Poly5_reg[56]  ( .D(n11470), .CP(clk), .CD(n18257), .Q(
        poly5_shifted[70]) );
  CFD2QXL \Poly5_reg[107]  ( .D(n11419), .CP(clk), .CD(n18260), .Q(
        poly5_shifted[121]) );
  CFD2QXL \Poly12_reg[69]  ( .D(n10463), .CP(clk), .CD(n18299), .Q(
        poly12_shifted[85]) );
  CFD2QXL \Poly1_reg[38]  ( .D(n9319), .CP(clk), .CD(n18373), .Q(
        poly1_shifted[49]) );
  CFD2QXL \polydata_reg[13]  ( .D(n8697), .CP(clk), .CD(n18257), .Q(
        polydata[13]) );
  CFD2QXL \polydata_reg[12]  ( .D(n8696), .CP(clk), .CD(n18257), .Q(
        polydata[12]) );
  CFD2QXL \Poly9_reg[98]  ( .D(n11207), .CP(clk), .CD(n18257), .Q(
        poly9_shifted[109]) );
  CFD2QXL \Poly12_reg[77]  ( .D(n10455), .CP(clk), .CD(n18297), .Q(
        poly12_shifted[93]) );
  CFD2QXL \Poly0_reg[126]  ( .D(n9451), .CP(clk), .CD(n18394), .Q(
        poly0_shifted[144]) );
  CFD2QXL \Poly0_reg[135]  ( .D(n9442), .CP(clk), .CD(n18394), .Q(
        poly0_shifted[153]) );
  CFD2QXL \Poly0_reg[37]  ( .D(n9540), .CP(clk), .CD(n18395), .Q(
        poly0_shifted[55]) );
  CFD2QXL \Poly0_reg[122]  ( .D(n9455), .CP(clk), .CD(n18394), .Q(
        poly0_shifted[140]) );
  CFD2QXL \Poly0_reg[144]  ( .D(n9433), .CP(clk), .CD(n18347), .Q(
        poly0_shifted[162]) );
  CFD2QXL \Poly1_reg[31]  ( .D(n9326), .CP(clk), .CD(n18368), .Q(
        poly1_shifted[42]) );
  CFD2QXL \Poly8_reg[37]  ( .D(n11364), .CP(clk), .CD(n18257), .Q(
        poly8_shifted[51]) );
  CFD2QXL \Poly3_reg[62]  ( .D(n8878), .CP(clk), .CD(n18381), .Q(
        poly3_shifted[76]) );
  CFD2QXL \Poly12_reg[48]  ( .D(n10484), .CP(clk), .CD(n18292), .Q(
        poly12_shifted[64]) );
  CFD2QXL \Poly14_reg[216]  ( .D(n10189), .CP(clk), .CD(n18303), .Q(
        poly14_shifted[232]) );
  CFD2QXL \Poly14_reg[230]  ( .D(n10175), .CP(clk), .CD(n18306), .Q(
        poly14_shifted[246]) );
  CFD2QXL \Poly13_reg[37]  ( .D(n11023), .CP(clk), .CD(n18281), .Q(
        poly13_shifted[51]) );
  CFD2QXL \Poly13_reg[51]  ( .D(n11009), .CP(clk), .CD(n18281), .Q(
        poly13_shifted[65]) );
  CFD2QXL \Poly13_reg[65]  ( .D(n10995), .CP(clk), .CD(n18281), .Q(
        poly13_shifted[79]) );
  CFD2QXL \Poly13_reg[79]  ( .D(n10981), .CP(clk), .CD(n18281), .Q(
        poly13_shifted[93]) );
  CFD2QXL \Poly13_reg[260]  ( .D(n10800), .CP(clk), .CD(n18286), .Q(
        poly13_shifted[274]) );
  CFD2QXL \Poly13_reg[5]  ( .D(n11055), .CP(clk), .CD(n18257), .Q(
        poly13_shifted[19]) );
  CFD2QXL \Poly13_reg[19]  ( .D(n11041), .CP(clk), .CD(n18257), .Q(
        poly13_shifted[33]) );
  CFD2QXL \Poly14_reg[11]  ( .D(n10394), .CP(clk), .CD(n18303), .Q(
        poly14_shifted[27]) );
  CFD2QXL \Poly14_reg[27]  ( .D(n10378), .CP(clk), .CD(n18303), .Q(
        poly14_shifted[43]) );
  CFD2QXL \Poly14_reg[43]  ( .D(n10362), .CP(clk), .CD(n18304), .Q(
        poly14_shifted[59]) );
  CFD2QXL \Poly14_reg[246]  ( .D(n10159), .CP(clk), .CD(n18306), .Q(
        poly14_shifted[262]) );
  CFD2QXL \Poly14_reg[262]  ( .D(n10143), .CP(clk), .CD(n18306), .Q(
        poly14_shifted[278]) );
  CFD2QXL \Poly14_reg[278]  ( .D(n10127), .CP(clk), .CD(n18306), .Q(
        poly14_shifted[294]) );
  CFD2QXL \Poly7_reg[132]  ( .D(n9972), .CP(clk), .CD(n18317), .Q(
        poly7_shifted[144]) );
  CFD2QXL \Poly7_reg[144]  ( .D(n9960), .CP(clk), .CD(n18317), .Q(
        poly7_shifted[156]) );
  CFD2QXL \Poly7_reg[156]  ( .D(n9948), .CP(clk), .CD(n18317), .Q(
        poly7_shifted[168]) );
  CFD2QXL \Poly7_reg[168]  ( .D(n9936), .CP(clk), .CD(n18317), .Q(
        poly7_shifted[180]) );
  CFD2QXL \Poly0_reg[0]  ( .D(n9577), .CP(clk), .CD(n18256), .Q(
        poly0_shifted[18]) );
  CFD2QXL \Poly0_reg[168]  ( .D(n9409), .CP(clk), .CD(n18348), .Q(
        poly0_shifted[186]) );
  CFD2QXL \Poly0_reg[4]  ( .D(n9573), .CP(clk), .CD(n18348), .Q(
        poly0_shifted[22]) );
  CFD2QXL \Poly0_reg[172]  ( .D(n9405), .CP(clk), .CD(n18348), .Q(
        poly0_shifted[190]) );
  CFD2QXL \Poly0_reg[169]  ( .D(n9408), .CP(clk), .CD(n18349), .Q(
        poly0_shifted[187]) );
  CFD2QXL \Poly0_reg[3]  ( .D(n9574), .CP(clk), .CD(n18349), .Q(
        poly0_shifted[21]) );
  CFD2QXL \Poly0_reg[147]  ( .D(n9430), .CP(clk), .CD(n18350), .Q(
        poly0_shifted[165]) );
  CFD2QXL \Poly0_reg[44]  ( .D(n9533), .CP(clk), .CD(n18350), .Q(
        poly0_shifted[62]) );
  CFD2QXL \Poly0_reg[171]  ( .D(n9406), .CP(clk), .CD(n18350), .Q(
        poly0_shifted[189]) );
  CFD2QXL \Poly0_reg[41]  ( .D(n9536), .CP(clk), .CD(n18350), .Q(
        poly0_shifted[59]) );
  CFD2QXL \Poly0_reg[149]  ( .D(n9428), .CP(clk), .CD(n18351), .Q(
        poly0_shifted[167]) );
  CFD2QXL \Poly0_reg[45]  ( .D(n9532), .CP(clk), .CD(n18352), .Q(
        poly0_shifted[63]) );
  CFD2QXL \Poly0_reg[142]  ( .D(n9435), .CP(clk), .CD(n18354), .Q(
        poly0_shifted[160]) );
  CFD2QXL \Poly0_reg[148]  ( .D(n9429), .CP(clk), .CD(n18357), .Q(
        poly0_shifted[166]) );
  CFD2QXL \Poly0_reg[1]  ( .D(n9576), .CP(clk), .CD(n18357), .Q(
        poly0_shifted[19]) );
  CFD2QXL \Poly0_reg[42]  ( .D(n9535), .CP(clk), .CD(n18357), .Q(
        poly0_shifted[60]) );
  CFD2QXL \Poly0_reg[140]  ( .D(n9437), .CP(clk), .CD(n18358), .Q(
        poly0_shifted[158]) );
  CFD2QXL \Poly0_reg[170]  ( .D(n9407), .CP(clk), .CD(n18348), .Q(
        poly0_shifted[188]) );
  CFD2QXL \dataselector_reg[34]  ( .D(n8761), .CP(clk), .CD(n18387), .Q(
        dataselector[34]) );
  CFD2QXL \dataselector_reg[48]  ( .D(n8747), .CP(clk), .CD(n18387), .Q(
        dataselector[48]) );
  CFD2QXL \dataselector_reg[32]  ( .D(n8763), .CP(clk), .CD(n18386), .Q(
        dataselector[32]) );
  CFD2QXL \dataselector_reg[10]  ( .D(n8785), .CP(clk), .CD(n18388), .Q(
        dataselector[10]) );
  CFD2QXL \dataselector_reg[46]  ( .D(n8749), .CP(clk), .CD(n18387), .Q(
        dataselector[46]) );
  CFD2QXL \Poly0_reg[174]  ( .D(n9403), .CP(clk), .CD(n18348), .Q(
        poly0_shifted[192]) );
  CFD2QXL \Poly0_reg[179]  ( .D(n9398), .CP(clk), .CD(n18393), .Q(
        poly0_shifted[197]) );
  CFD2QXL \Poly10_reg[23]  ( .D(n11080), .CP(clk), .CD(n18262), .Q(Poly10[23])
         );
  CFD2QXL \Poly13_reg[2]  ( .D(n11058), .CP(clk), .CD(n18269), .Q(
        poly13_shifted[16]) );
  CFD2QXL \Poly14_reg[23]  ( .D(n10382), .CP(clk), .CD(n18301), .Q(
        poly14_shifted[39]) );
  CFD2QXL \Poly12_reg[119]  ( .D(n10413), .CP(clk), .CD(n18295), .Q(
        Poly12[119]) );
  CFD2QXL \Poly2_reg[49]  ( .D(n8961), .CP(clk), .CD(n18379), .Q(Poly2[49]) );
  CFD2QXL \dataselector_reg[50]  ( .D(n8745), .CP(clk), .CD(n18257), .Q(
        dataselector[50]) );
  CFD2QXL \dataselector_reg[55]  ( .D(n8740), .CP(clk), .CD(n18257), .Q(
        dataselector[55]) );
  CFD2QXL \polydata_reg[11]  ( .D(n8695), .CP(clk), .CD(n18401), .Q(
        polydata[11]) );
  CFD2QXL \polydata_reg[2]  ( .D(n8686), .CP(clk), .CD(n18401), .Q(polydata[2]) );
  CFD2QXL \Poly11_reg[75]  ( .D(n11114), .CP(clk), .CD(n18257), .Q(Poly11[75])
         );
  CFD2QXL \Poly10_reg[9]  ( .D(n11094), .CP(clk), .CD(n18263), .Q(
        poly10_shifted[21]) );
  CFD2QXL \Poly2_reg[61]  ( .D(n8949), .CP(clk), .CD(n18380), .Q(Poly2[61]) );
  CFD2QXL \Poly4_reg[36]  ( .D(n8820), .CP(clk), .CD(n18389), .Q(Poly4[36]) );
  CFD2QXL \dataselector_reg[19]  ( .D(n8776), .CP(clk), .CD(n18388), .Q(
        dataselector[19]) );
  CFD2QXL \Poly10_reg[32]  ( .D(n11071), .CP(clk), .CD(n18262), .Q(Poly10[32])
         );
  CFD2QXL \Poly5_reg[31]  ( .D(n11495), .CP(clk), .CD(n18257), .Q(
        poly5_shifted[45]) );
  CFD2QXL \Poly5_reg[52]  ( .D(n11474), .CP(clk), .CD(n18260), .Q(
        poly5_shifted[66]) );
  CFD2QXL \Poly10_reg[20]  ( .D(n11083), .CP(clk), .CD(n18263), .Q(Poly10[20])
         );
  CFD2QXL \Poly7_reg[349]  ( .D(n9755), .CP(clk), .CD(n18336), .Q(
        poly7_shifted[361]) );
  CFD2QXL \Poly15_reg[15]  ( .D(n9622), .CP(clk), .CD(n18344), .Q(Poly15[15])
         );
  CFD2QXL \Poly0_reg[71]  ( .D(n9506), .CP(clk), .CD(n18356), .Q(
        poly0_shifted[89]) );
  CFD2QXL \Poly5_reg[101]  ( .D(n11425), .CP(clk), .CD(n18257), .Q(Poly5[101])
         );
  CFD2QXL \Poly5_reg[102]  ( .D(n11424), .CP(clk), .CD(n18257), .Q(Poly5[102])
         );
  CFD2QXL \Poly8_reg[16]  ( .D(n11385), .CP(clk), .CD(n18257), .Q(Poly8[16])
         );
  CFD2QXL \Poly9_reg[25]  ( .D(n11280), .CP(clk), .CD(n18257), .Q(Poly9[25])
         );
  CFD2QXL \Poly9_reg[26]  ( .D(n11279), .CP(clk), .CD(n18257), .Q(Poly9[26])
         );
  CFD2QXL \Poly11_reg[66]  ( .D(n11123), .CP(clk), .CD(n18257), .Q(Poly11[66])
         );
  CFD2QXL \Poly10_reg[24]  ( .D(n11079), .CP(clk), .CD(n18400), .Q(Poly10[24])
         );
  CFD2QXL \Poly10_reg[21]  ( .D(n11082), .CP(clk), .CD(n18263), .Q(Poly10[21])
         );
  CFD2QXL \Poly10_reg[26]  ( .D(n11077), .CP(clk), .CD(n18263), .Q(Poly10[26])
         );
  CFD2QXL \Poly10_reg[19]  ( .D(n11084), .CP(clk), .CD(n18263), .Q(Poly10[19])
         );
  CFD2QXL \Poly12_reg[35]  ( .D(n10497), .CP(clk), .CD(n18294), .Q(Poly12[35])
         );
  CFD2QXL \Poly12_reg[67]  ( .D(n10465), .CP(clk), .CD(n18298), .Q(Poly12[67])
         );
  CFD2QXL \Poly14_reg[195]  ( .D(n10210), .CP(clk), .CD(n18314), .Q(
        Poly14[195]) );
  CFD2QXL \Poly6_reg[36]  ( .D(n9657), .CP(clk), .CD(n18344), .Q(Poly6[36]) );
  CFD2QXL \Poly2_reg[35]  ( .D(n8975), .CP(clk), .CD(n18380), .Q(Poly2[35]) );
  CFD2QXL \Poly3_reg[48]  ( .D(n8892), .CP(clk), .CD(n18381), .Q(Poly3[48]) );
  CFD2QXL \Poly5_reg[19]  ( .D(n11507), .CP(clk), .CD(n18257), .Q(
        poly5_shifted[33]) );
  CFD2QXL \Poly5_reg[26]  ( .D(n11500), .CP(clk), .CD(n18257), .Q(
        poly5_shifted[40]) );
  CFD2QXL \Poly0_reg[101]  ( .D(n9476), .CP(clk), .CD(n18394), .Q(
        poly0_shifted[119]) );
  CFD2QXL \Poly0_reg[69]  ( .D(n9508), .CP(clk), .CD(n18355), .Q(
        poly0_shifted[87]) );
  CFD2QXL \Poly2_reg[16]  ( .D(n8994), .CP(clk), .CD(n18378), .Q(
        poly2_shifted[28]) );
  CFD2QXL \Poly6_reg[35]  ( .D(n9658), .CP(clk), .CD(n18344), .Q(Poly6[35]) );
  CFD2QXL \dataselector_reg[36]  ( .D(n8759), .CP(clk), .CD(n18387), .Q(
        dataselector[36]) );
  CFD2QXL \Poly12_reg[41]  ( .D(n10491), .CP(clk), .CD(n18296), .Q(
        poly12_shifted[57]) );
  CFD2QXL \Poly7_reg[315]  ( .D(n9789), .CP(clk), .CD(n18339), .Q(
        poly7_shifted[327]) );
  CFD2QXL \Poly2_reg[57]  ( .D(n8953), .CP(clk), .CD(n18379), .Q(Poly2[57]) );
  CFD2QXL \Poly2_reg[28]  ( .D(n8982), .CP(clk), .CD(n18391), .Q(Poly2[28]) );
  CFD2QXL \Poly0_reg[180]  ( .D(n9397), .CP(clk), .CD(n18347), .Q(
        poly0_shifted[198]) );
  CFD2QXL \dataselector_reg[0]  ( .D(n8795), .CP(clk), .CD(n18386), .Q(
        dataselector[0]) );
  CFD2QXL \Poly0_reg[208]  ( .D(n9369), .CP(clk), .CD(n18348), .Q(Poly0[208])
         );
  CFD2QXL \dataselector_reg[15]  ( .D(n8780), .CP(clk), .CD(n18388), .Q(
        dataselector[15]) );
  CFD2QXL \dataselector_reg[4]  ( .D(n8791), .CP(clk), .CD(n18386), .Q(
        dataselector[4]) );
  CFD2QXL \dataselector_reg[24]  ( .D(n8771), .CP(clk), .CD(n18387), .Q(
        dataselector[24]) );
  CFD2QXL \dataselector_reg[27]  ( .D(n8768), .CP(clk), .CD(n18387), .Q(
        dataselector[27]) );
  CFD2QXL \Poly5_reg[70]  ( .D(n11456), .CP(clk), .CD(n18257), .Q(
        poly5_shifted[84]) );
  CFD2QXL \Poly5_reg[33]  ( .D(n11493), .CP(clk), .CD(n18257), .Q(
        poly5_shifted[47]) );
  CFD2QXL \Poly5_reg[103]  ( .D(n11423), .CP(clk), .CD(n18257), .Q(
        poly5_shifted[117]) );
  CFD2QXL \Poly5_reg[40]  ( .D(n11486), .CP(clk), .CD(n18257), .Q(
        poly5_shifted[54]) );
  CFD2QXL \Poly5_reg[66]  ( .D(n11460), .CP(clk), .CD(n18260), .Q(
        poly5_shifted[80]) );
  CFD2QXL \Poly6_reg[37]  ( .D(n9656), .CP(clk), .CD(n18343), .Q(Poly6[37]) );
  CFD2QXL \Poly2_reg[52]  ( .D(n8958), .CP(clk), .CD(n18378), .Q(Poly2[52]) );
  CFD2QXL \Poly2_reg[53]  ( .D(n8957), .CP(clk), .CD(n18380), .Q(Poly2[53]) );
  CFD2QXL \Poly2_reg[51]  ( .D(n8959), .CP(clk), .CD(n18380), .Q(Poly2[51]) );
  CFD2QXL \Poly4_reg[43]  ( .D(n8813), .CP(clk), .CD(n18385), .Q(Poly4[43]) );
  CFD2QXL \dataselector_reg[28]  ( .D(n8767), .CP(clk), .CD(n18388), .Q(
        dataselector[28]) );
  CFD2QXL \scrambler_reg[1]  ( .D(n8701), .CP(clk), .CD(n18257), .Q(
        scrambler[1]) );
  CFD2QXL \Poly11_reg[55]  ( .D(n11134), .CP(clk), .CD(n18257), .Q(Poly11[55])
         );
  CFD2QXL \Poly2_reg[33]  ( .D(n8977), .CP(clk), .CD(n18379), .Q(Poly2[33]) );
  CFD2QXL \Poly3_reg[45]  ( .D(n8895), .CP(clk), .CD(n18381), .Q(Poly3[45]) );
  CFD2QXL \Poly3_reg[47]  ( .D(n8893), .CP(clk), .CD(n18384), .Q(Poly3[47]) );
  CFD2QXL \Poly3_reg[50]  ( .D(n8890), .CP(clk), .CD(n18384), .Q(Poly3[50]) );
  CFD2QXL \Poly4_reg[42]  ( .D(n8814), .CP(clk), .CD(n18385), .Q(Poly4[42]) );
  CFD2QXL \Poly2_reg[55]  ( .D(n8955), .CP(clk), .CD(n18379), .Q(Poly2[55]) );
  CFD2QXL \Poly0_reg[191]  ( .D(n9386), .CP(clk), .CD(n18393), .Q(
        poly0_shifted[209]) );
  CFD2QXL \Poly0_reg[63]  ( .D(n9514), .CP(clk), .CD(n18394), .Q(
        poly0_shifted[81]) );
  CFD2QXL \dataselector_reg[33]  ( .D(n8762), .CP(clk), .CD(n18388), .Q(
        dataselector[33]) );
  CFD2QXL \scrambler_reg[11]  ( .D(n8711), .CP(clk), .CD(n18401), .Q(
        scrambler[11]) );
  CFD2QXL \Poly0_reg[165]  ( .D(n9412), .CP(clk), .CD(n18350), .Q(Poly0[165])
         );
  CFD2QXL \Poly0_reg[19]  ( .D(n9558), .CP(clk), .CD(n18357), .Q(Poly0[19]) );
  CFD2QXL \Poly0_reg[54]  ( .D(n9523), .CP(clk), .CD(n18395), .Q(
        poly0_shifted[72]) );
  CFD2QXL \Poly0_reg[186]  ( .D(n9391), .CP(clk), .CD(n18394), .Q(
        poly0_shifted[204]) );
  CFD2QXL \Poly0_reg[188]  ( .D(n9389), .CP(clk), .CD(n18394), .Q(
        poly0_shifted[206]) );
  CFD2QXL \Poly0_reg[187]  ( .D(n9390), .CP(clk), .CD(n18394), .Q(
        poly0_shifted[205]) );
  CFD2QXL \Poly0_reg[57]  ( .D(n9520), .CP(clk), .CD(n18395), .Q(
        poly0_shifted[75]) );
  CFD2QXL \Poly0_reg[62]  ( .D(n9515), .CP(clk), .CD(n18394), .Q(
        poly0_shifted[80]) );
  CFD2QXL \Poly0_reg[189]  ( .D(n9388), .CP(clk), .CD(n18394), .Q(
        poly0_shifted[207]) );
  CFD2QXL \Poly0_reg[59]  ( .D(n9518), .CP(clk), .CD(n18395), .Q(
        poly0_shifted[77]) );
  CFD2QXL \Poly0_reg[61]  ( .D(n9516), .CP(clk), .CD(n18394), .Q(
        poly0_shifted[79]) );
  CFD2QXL \Poly0_reg[48]  ( .D(n9529), .CP(clk), .CD(n18395), .Q(
        poly0_shifted[66]) );
  CFD2QXL \Poly0_reg[47]  ( .D(n9530), .CP(clk), .CD(n18395), .Q(
        poly0_shifted[65]) );
  CFD2QXL \Poly0_reg[49]  ( .D(n9528), .CP(clk), .CD(n18395), .Q(
        poly0_shifted[67]) );
  CFD2QXL \Poly0_reg[51]  ( .D(n9526), .CP(clk), .CD(n18395), .Q(
        poly0_shifted[69]) );
  CFD2QXL \Poly0_reg[56]  ( .D(n9521), .CP(clk), .CD(n18395), .Q(
        poly0_shifted[74]) );
  CFD2QXL \Poly0_reg[53]  ( .D(n9524), .CP(clk), .CD(n18395), .Q(
        poly0_shifted[71]) );
  CFD2QXL \Poly0_reg[58]  ( .D(n9519), .CP(clk), .CD(n18395), .Q(
        poly0_shifted[76]) );
  CFD2QXL \Poly0_reg[55]  ( .D(n9522), .CP(clk), .CD(n18395), .Q(
        poly0_shifted[73]) );
  CFD2QXL \Poly0_reg[60]  ( .D(n9517), .CP(clk), .CD(n18395), .Q(
        poly0_shifted[78]) );
  CFD2QXL \Poly8_reg[43]  ( .D(n11358), .CP(clk), .CD(n18257), .Q(
        poly8_shifted[57]) );
  CFD2QXL \Poly13_reg[14]  ( .D(n11046), .CP(clk), .CD(n18264), .Q(
        poly13_shifted[28]) );
  CFD2QXL \Poly13_reg[18]  ( .D(n11042), .CP(clk), .CD(n18266), .Q(
        poly13_shifted[32]) );
  CFD2QXL \Poly13_reg[29]  ( .D(n11031), .CP(clk), .CD(n18270), .Q(
        poly13_shifted[43]) );
  CFD2QXL \Poly13_reg[27]  ( .D(n11033), .CP(clk), .CD(n18274), .Q(
        poly13_shifted[41]) );
  CFD2QXL \Poly12_reg[76]  ( .D(n10456), .CP(clk), .CD(n18296), .Q(
        poly12_shifted[92]) );
  CFD2QXL \Poly7_reg[303]  ( .D(n9801), .CP(clk), .CD(n18339), .Q(
        poly7_shifted[315]) );
  CFD2QXL \Poly7_reg[43]  ( .D(n10061), .CP(clk), .CD(n18340), .Q(
        poly7_shifted[55]) );
  CFD2QXL \Poly7_reg[103]  ( .D(n10001), .CP(clk), .CD(n18340), .Q(
        poly7_shifted[115]) );
  CFD2QXL \Poly1_reg[44]  ( .D(n9313), .CP(clk), .CD(n18358), .Q(
        poly1_shifted[55]) );
  CFD2QXL \Poly1_reg[279]  ( .D(n9078), .CP(clk), .CD(n18367), .Q(
        poly1_shifted[290]) );
  CFD2QXL \Poly1_reg[256]  ( .D(n9101), .CP(clk), .CD(n18369), .Q(
        poly1_shifted[267]) );
  CFD2QXL \Poly1_reg[289]  ( .D(n9068), .CP(clk), .CD(n18369), .Q(
        poly1_shifted[300]) );
  CFD2QXL \Poly0_reg[175]  ( .D(n9402), .CP(clk), .CD(n18393), .Q(
        poly0_shifted[193]) );
  CFD2QXL \Poly0_reg[157]  ( .D(n9420), .CP(clk), .CD(n18354), .Q(Poly0[157])
         );
  CFD2QXL \dataselector_reg[26]  ( .D(n8769), .CP(clk), .CD(n18386), .Q(
        dataselector[26]) );
  CFD2QXL \dataselector_reg[2]  ( .D(n8793), .CP(clk), .CD(n18388), .Q(
        dataselector[2]) );
  CFD2QXL \dataselector_reg[23]  ( .D(n8772), .CP(clk), .CD(n18387), .Q(
        dataselector[23]) );
  CFD2QXL \dataselector_reg[6]  ( .D(n8789), .CP(clk), .CD(n18387), .Q(
        dataselector[6]) );
  CFD2QXL \Poly7_reg[339]  ( .D(n9765), .CP(clk), .CD(n18339), .Q(
        poly7_shifted[351]) );
  CFD2QXL \Poly5_reg[63]  ( .D(n11463), .CP(clk), .CD(n18257), .Q(
        poly5_shifted[77]) );
  CFD2QXL \Poly5_reg[6]  ( .D(n11520), .CP(clk), .CD(n18257), .Q(
        poly5_shifted[20]) );
  CFD2QXL \Poly7_reg[361]  ( .D(n9743), .CP(clk), .CD(n18336), .Q(
        poly7_shifted[373]) );
  CFD2QXL \Poly0_reg[89]  ( .D(n9488), .CP(clk), .CD(n18356), .Q(
        poly0_shifted[107]) );
  CFD2QXL \Poly0_reg[182]  ( .D(n9395), .CP(clk), .CD(n18347), .Q(
        poly0_shifted[200]) );
  CFD2QXL \Poly0_reg[177]  ( .D(n9400), .CP(clk), .CD(n18353), .Q(
        poly0_shifted[195]) );
  CFD2QXL \Poly0_reg[185]  ( .D(n9392), .CP(clk), .CD(n18357), .Q(
        poly0_shifted[203]) );
  CFD2QXL \Poly8_reg[32]  ( .D(n11369), .CP(clk), .CD(n18257), .Q(
        poly8_shifted[46]) );
  CFD2QXL \Poly7_reg[31]  ( .D(n10073), .CP(clk), .CD(n18339), .Q(
        poly7_shifted[43]) );
  CFD2QXL \Poly13_reg[49]  ( .D(n11011), .CP(clk), .CD(n18285), .Q(
        poly13_shifted[63]) );
  CFD2QXL \Poly14_reg[15]  ( .D(n10390), .CP(clk), .CD(n18305), .Q(
        poly14_shifted[31]) );
  CFD2QXL \Poly0_reg[43]  ( .D(n9534), .CP(clk), .CD(n18351), .Q(
        poly0_shifted[61]) );
  CFD2QXL \Poly0_reg[124]  ( .D(n9453), .CP(clk), .CD(n18354), .Q(
        poly0_shifted[142]) );
  CFD2QXL \Poly0_reg[121]  ( .D(n9456), .CP(clk), .CD(n18354), .Q(
        poly0_shifted[139]) );
  CFD2QXL \Poly0_reg[141]  ( .D(n9436), .CP(clk), .CD(n18355), .Q(
        poly0_shifted[159]) );
  CFD2QXL \Poly3_reg[59]  ( .D(n8881), .CP(clk), .CD(n18380), .Q(
        poly3_shifted[73]) );
  CFD2QXL \Poly13_reg[468]  ( .D(n10592), .CP(clk), .CD(n18278), .Q(
        poly13_shifted[482]) );
  CFD2QXL \Poly13_reg[23]  ( .D(n11037), .CP(clk), .CD(n18281), .Q(
        poly13_shifted[37]) );
  CFD2QXL \Poly13_reg[246]  ( .D(n10814), .CP(clk), .CD(n18285), .Q(
        poly13_shifted[260]) );
  CFD2QXL \Poly13_reg[505]  ( .D(n10555), .CP(clk), .CD(n18289), .Q(
        poly13_shifted[519]) );
  CFD2QXL \Poly14_reg[161]  ( .D(n10244), .CP(clk), .CD(n18303), .Q(
        poly14_shifted[177]) );
  CFD2QXL \Poly14_reg[280]  ( .D(n10125), .CP(clk), .CD(n18303), .Q(
        poly14_shifted[296]) );
  CFD2QXL \Poly14_reg[159]  ( .D(n10246), .CP(clk), .CD(n18306), .Q(
        poly14_shifted[175]) );
  CFD2QXL \Poly7_reg[120]  ( .D(n9984), .CP(clk), .CD(n18317), .Q(
        poly7_shifted[132]) );
  CFD2QXL \Poly2_reg[45]  ( .D(n8965), .CP(clk), .CD(n18379), .Q(
        poly2_shifted[57]) );
  CFD2QXL \Poly5_reg[90]  ( .D(n11436), .CP(clk), .CD(n18257), .Q(Poly5[90])
         );
  CFD2QXL \Poly5_reg[110]  ( .D(n11416), .CP(clk), .CD(n18257), .Q(
        poly5_shifted[124]) );
  CFD2QXL \Poly5_reg[108]  ( .D(n11418), .CP(clk), .CD(n18258), .Q(
        poly5_shifted[122]) );
  CFD2QXL \Poly5_reg[106]  ( .D(n11420), .CP(clk), .CD(n18258), .Q(
        poly5_shifted[120]) );
  CFD2QXL \Poly5_reg[17]  ( .D(n11509), .CP(clk), .CD(n18257), .Q(
        poly5_shifted[31]) );
  CFD2QXL \Poly5_reg[18]  ( .D(n11508), .CP(clk), .CD(n18257), .Q(
        poly5_shifted[32]) );
  CFD2QXL \Poly8_reg[0]  ( .D(n11401), .CP(clk), .CD(n18257), .Q(
        poly8_shifted[14]) );
  CFD2QXL \Poly8_reg[28]  ( .D(n11373), .CP(clk), .CD(n18257), .Q(
        poly8_shifted[42]) );
  CFD2QXL \Poly8_reg[26]  ( .D(n11375), .CP(clk), .CD(n18261), .Q(
        poly8_shifted[40]) );
  CFD2QXL \Poly9_reg[99]  ( .D(n11206), .CP(clk), .CD(n18257), .Q(
        poly9_shifted[110]) );
  CFD2QXL \Poly9_reg[32]  ( .D(n11273), .CP(clk), .CD(n18257), .Q(
        poly9_shifted[43]) );
  CFD2QXL \Poly9_reg[95]  ( .D(n11210), .CP(clk), .CD(n18257), .Q(
        poly9_shifted[106]) );
  CFD2QXL \Poly9_reg[34]  ( .D(n11271), .CP(clk), .CD(n18257), .Q(
        poly9_shifted[45]) );
  CFD2QXL \Poly9_reg[96]  ( .D(n11209), .CP(clk), .CD(n18257), .Q(
        poly9_shifted[107]) );
  CFD2QXL \Poly10_reg[29]  ( .D(n11074), .CP(clk), .CD(n18263), .Q(
        poly10_shifted[41]) );
  CFD2QXL \Poly13_reg[182]  ( .D(n10878), .CP(clk), .CD(n18265), .Q(
        poly13_shifted[196]) );
  CFD2QXL \Poly13_reg[406]  ( .D(n10654), .CP(clk), .CD(n18266), .Q(
        poly13_shifted[420]) );
  CFD2QXL \Poly13_reg[172]  ( .D(n10888), .CP(clk), .CD(n18268), .Q(
        poly13_shifted[186]) );
  CFD2QXL \Poly13_reg[171]  ( .D(n10889), .CP(clk), .CD(n18257), .Q(
        poly13_shifted[185]) );
  CFD2QXL \Poly13_reg[284]  ( .D(n10776), .CP(clk), .CD(n18271), .Q(
        poly13_shifted[298]) );
  CFD2QXL \Poly13_reg[402]  ( .D(n10658), .CP(clk), .CD(n18272), .Q(
        poly13_shifted[416]) );
  CFD2QXL \Poly13_reg[169]  ( .D(n10891), .CP(clk), .CD(n18272), .Q(
        poly13_shifted[183]) );
  CFD2QXL \Poly13_reg[401]  ( .D(n10659), .CP(clk), .CD(n18273), .Q(
        poly13_shifted[415]) );
  CFD2QXL \Poly13_reg[296]  ( .D(n10764), .CP(clk), .CD(n18275), .Q(
        poly13_shifted[310]) );
  CFD2QXL \Poly13_reg[295]  ( .D(n10765), .CP(clk), .CD(n18255), .Q(
        poly13_shifted[309]) );
  CFD2QXL \Poly13_reg[412]  ( .D(n10648), .CP(clk), .CD(n18278), .Q(
        poly13_shifted[426]) );
  CFD2QXL \Poly13_reg[178]  ( .D(n10882), .CP(clk), .CD(n18282), .Q(
        poly13_shifted[192]) );
  CFD2QXL \Poly13_reg[410]  ( .D(n10650), .CP(clk), .CD(n18283), .Q(
        poly13_shifted[424]) );
  CFD2QXL \Poly13_reg[177]  ( .D(n10883), .CP(clk), .CD(n18255), .Q(
        poly13_shifted[191]) );
  CFD2QXL \Poly13_reg[291]  ( .D(n10769), .CP(clk), .CD(n18255), .Q(
        poly13_shifted[305]) );
  CFD2QXL \Poly13_reg[176]  ( .D(n10884), .CP(clk), .CD(n18285), .Q(
        poly13_shifted[190]) );
  CFD2QXL \Poly13_reg[290]  ( .D(n10770), .CP(clk), .CD(n18286), .Q(
        poly13_shifted[304]) );
  CFD2QXL \Poly13_reg[175]  ( .D(n10885), .CP(clk), .CD(n18287), .Q(
        poly13_shifted[189]) );
  CFD2QXL \Poly13_reg[287]  ( .D(n10773), .CP(clk), .CD(n18288), .Q(
        poly13_shifted[301]) );
  CFD2QXL \Poly13_reg[407]  ( .D(n10653), .CP(clk), .CD(n18289), .Q(
        poly13_shifted[421]) );
  CFD2QXL \Poly13_reg[288]  ( .D(n10772), .CP(clk), .CD(n18291), .Q(
        poly13_shifted[302]) );
  CFD2QXL \Poly12_reg[80]  ( .D(n10452), .CP(clk), .CD(n18292), .Q(
        poly12_shifted[96]) );
  CFD2QXL \Poly12_reg[9]  ( .D(n10523), .CP(clk), .CD(n18293), .Q(
        poly12_shifted[25]) );
  CFD2QXL \Poly12_reg[11]  ( .D(n10521), .CP(clk), .CD(n18293), .Q(
        poly12_shifted[27]) );
  CFD2QXL \Poly12_reg[12]  ( .D(n10520), .CP(clk), .CD(n18296), .Q(
        poly12_shifted[28]) );
  CFD2QXL \Poly12_reg[44]  ( .D(n10488), .CP(clk), .CD(n18296), .Q(
        poly12_shifted[60]) );
  CFD2QXL \Poly12_reg[78]  ( .D(n10454), .CP(clk), .CD(n18297), .Q(
        poly12_shifted[94]) );
  CFD2QXL \Poly12_reg[45]  ( .D(n10487), .CP(clk), .CD(n18297), .Q(
        poly12_shifted[61]) );
  CFD2QXL \Poly12_reg[79]  ( .D(n10453), .CP(clk), .CD(n18298), .Q(
        poly12_shifted[95]) );
  CFD2QXL \Poly12_reg[2]  ( .D(n10530), .CP(clk), .CD(n18298), .Q(
        poly12_shifted[18]) );
  CFD2QXL \Poly12_reg[50]  ( .D(n10482), .CP(clk), .CD(n18298), .Q(
        poly12_shifted[66]) );
  CFD2QXL \Poly12_reg[49]  ( .D(n10483), .CP(clk), .CD(n18298), .Q(
        poly12_shifted[65]) );
  CFD2QXL \Poly12_reg[40]  ( .D(n10492), .CP(clk), .CD(n18299), .Q(
        poly12_shifted[56]) );
  CFD2QXL \Poly12_reg[70]  ( .D(n10462), .CP(clk), .CD(n18299), .Q(
        poly12_shifted[86]) );
  CFD2QXL \Poly14_reg[7]  ( .D(n10398), .CP(clk), .CD(n18301), .Q(
        poly14_shifted[23]) );
  CFD2QXL \Poly14_reg[222]  ( .D(n10183), .CP(clk), .CD(n18302), .Q(
        poly14_shifted[238]) );
  CFD2QXL \Poly14_reg[1]  ( .D(n10404), .CP(clk), .CD(n18302), .Q(
        poly14_shifted[17]) );
  CFD2QXL \Poly14_reg[5]  ( .D(n10400), .CP(clk), .CD(n18304), .Q(
        poly14_shifted[21]) );
  CFD2QXL \Poly14_reg[220]  ( .D(n10185), .CP(clk), .CD(n18305), .Q(
        poly14_shifted[236]) );
  CFD2QXL \Poly14_reg[185]  ( .D(n10220), .CP(clk), .CD(n18307), .Q(
        poly14_shifted[201]) );
  CFD2QXL \Poly14_reg[217]  ( .D(n10188), .CP(clk), .CD(n18307), .Q(
        poly14_shifted[233]) );
  CFD2QXL \Poly14_reg[188]  ( .D(n10217), .CP(clk), .CD(n18308), .Q(
        poly14_shifted[204]) );
  CFD2QXL \Poly14_reg[227]  ( .D(n10178), .CP(clk), .CD(n18308), .Q(
        poly14_shifted[243]) );
  CFD2QXL \Poly14_reg[182]  ( .D(n10223), .CP(clk), .CD(n18309), .Q(
        poly14_shifted[198]) );
  CFD2QXL \Poly14_reg[186]  ( .D(n10219), .CP(clk), .CD(n18311), .Q(
        poly14_shifted[202]) );
  CFD2QXL \Poly14_reg[191]  ( .D(n10214), .CP(clk), .CD(n18311), .Q(
        poly14_shifted[207]) );
  CFD2QXL \Poly14_reg[225]  ( .D(n10180), .CP(clk), .CD(n18311), .Q(
        poly14_shifted[241]) );
  CFD2QXL \Poly14_reg[229]  ( .D(n10176), .CP(clk), .CD(n18314), .Q(
        poly14_shifted[245]) );
  CFD2QXL \Poly14_reg[8]  ( .D(n10397), .CP(clk), .CD(n18314), .Q(
        poly14_shifted[24]) );
  CFD2QXL \Poly14_reg[223]  ( .D(n10182), .CP(clk), .CD(n18315), .Q(
        poly14_shifted[239]) );
  CFD2QXL \Poly14_reg[183]  ( .D(n10222), .CP(clk), .CD(n18316), .Q(
        poly14_shifted[199]) );
  CFD2QXL \Poly7_reg[36]  ( .D(n10068), .CP(clk), .CD(n18316), .Q(
        poly7_shifted[48]) );
  CFD2QXL \Poly7_reg[60]  ( .D(n10044), .CP(clk), .CD(n18317), .Q(
        poly7_shifted[72]) );
  CFD2QXL \Poly7_reg[204]  ( .D(n9900), .CP(clk), .CD(n18317), .Q(
        poly7_shifted[216]) );
  CFD2QXL \Poly7_reg[252]  ( .D(n9852), .CP(clk), .CD(n18318), .Q(
        poly7_shifted[264]) );
  CFD2QXL \Poly7_reg[254]  ( .D(n9850), .CP(clk), .CD(n18319), .Q(
        poly7_shifted[266]) );
  CFD2QXL \Poly7_reg[11]  ( .D(n10093), .CP(clk), .CD(n18319), .Q(
        poly7_shifted[23]) );
  CFD2QXL \Poly7_reg[256]  ( .D(n9848), .CP(clk), .CD(n18319), .Q(
        poly7_shifted[268]) );
  CFD2QXL \Poly7_reg[246]  ( .D(n9858), .CP(clk), .CD(n18320), .Q(
        poly7_shifted[258]) );
  CFD2QXL \Poly7_reg[248]  ( .D(n9856), .CP(clk), .CD(n18321), .Q(
        poly7_shifted[260]) );
  CFD2QXL \Poly7_reg[5]  ( .D(n10099), .CP(clk), .CD(n18322), .Q(
        poly7_shifted[17]) );
  CFD2QXL \Poly7_reg[250]  ( .D(n9854), .CP(clk), .CD(n18322), .Q(
        poly7_shifted[262]) );
  CFD2QXL \Poly7_reg[38]  ( .D(n10066), .CP(clk), .CD(n18325), .Q(
        poly7_shifted[50]) );
  CFD2QXL \Poly7_reg[33]  ( .D(n10071), .CP(clk), .CD(n18325), .Q(
        poly7_shifted[45]) );
  CFD2QXL \Poly7_reg[69]  ( .D(n10035), .CP(clk), .CD(n18325), .Q(
        poly7_shifted[81]) );
  CFD2QXL \Poly7_reg[62]  ( .D(n10042), .CP(clk), .CD(n18326), .Q(
        poly7_shifted[74]) );
  CFD2QXL \Poly7_reg[247]  ( .D(n9857), .CP(clk), .CD(n18326), .Q(
        poly7_shifted[259]) );
  CFD2QXL \Poly7_reg[35]  ( .D(n10069), .CP(clk), .CD(n18328), .Q(
        poly7_shifted[47]) );
  CFD2QXL \Poly7_reg[71]  ( .D(n10033), .CP(clk), .CD(n18328), .Q(
        poly7_shifted[83]) );
  CFD2QXL \Poly7_reg[64]  ( .D(n10040), .CP(clk), .CD(n18328), .Q(
        poly7_shifted[76]) );
  CFD2QXL \Poly7_reg[206]  ( .D(n9898), .CP(clk), .CD(n18329), .Q(
        poly7_shifted[218]) );
  CFD2QXL \Poly7_reg[249]  ( .D(n9855), .CP(clk), .CD(n18329), .Q(
        poly7_shifted[261]) );
  CFD2QXL \Poly7_reg[42]  ( .D(n10062), .CP(clk), .CD(n18330), .Q(
        poly7_shifted[54]) );
  CFD2QXL \Poly7_reg[37]  ( .D(n10067), .CP(clk), .CD(n18331), .Q(
        poly7_shifted[49]) );
  CFD2QXL \Poly7_reg[66]  ( .D(n10038), .CP(clk), .CD(n18331), .Q(
        poly7_shifted[78]) );
  CFD2QXL \Poly7_reg[196]  ( .D(n9908), .CP(clk), .CD(n18332), .Q(
        poly7_shifted[208]) );
  CFD2QXL \Poly7_reg[201]  ( .D(n9903), .CP(clk), .CD(n18332), .Q(
        poly7_shifted[213]) );
  CFD2QXL \Poly7_reg[32]  ( .D(n10072), .CP(clk), .CD(n18334), .Q(
        poly7_shifted[44]) );
  CFD2QXL \Poly7_reg[39]  ( .D(n10065), .CP(clk), .CD(n18334), .Q(
        poly7_shifted[51]) );
  CFD2QXL \Poly7_reg[63]  ( .D(n10041), .CP(clk), .CD(n18334), .Q(
        poly7_shifted[75]) );
  CFD2QXL \Poly7_reg[68]  ( .D(n10036), .CP(clk), .CD(n18335), .Q(
        poly7_shifted[80]) );
  CFD2QXL \Poly7_reg[203]  ( .D(n9901), .CP(clk), .CD(n18335), .Q(
        poly7_shifted[215]) );
  CFD2QXL \Poly7_reg[34]  ( .D(n10070), .CP(clk), .CD(n18337), .Q(
        poly7_shifted[46]) );
  CFD2QXL \Poly7_reg[41]  ( .D(n10063), .CP(clk), .CD(n18337), .Q(
        poly7_shifted[53]) );
  CFD2QXL \Poly7_reg[65]  ( .D(n10039), .CP(clk), .CD(n18337), .Q(
        poly7_shifted[77]) );
  CFD2QXL \Poly7_reg[70]  ( .D(n10034), .CP(clk), .CD(n18338), .Q(
        poly7_shifted[82]) );
  CFD2QXL \Poly7_reg[200]  ( .D(n9904), .CP(clk), .CD(n18338), .Q(
        poly7_shifted[212]) );
  CFD2QXL \Poly7_reg[205]  ( .D(n9899), .CP(clk), .CD(n18338), .Q(
        poly7_shifted[217]) );
  CFD2QXL \Poly7_reg[255]  ( .D(n9849), .CP(clk), .CD(n18339), .Q(
        poly7_shifted[267]) );
  CFD2QXL \Poly7_reg[195]  ( .D(n9909), .CP(clk), .CD(n18341), .Q(
        poly7_shifted[207]) );
  CFD2QXL \Poly7_reg[202]  ( .D(n9902), .CP(clk), .CD(n18341), .Q(
        poly7_shifted[214]) );
  CFD2QXL \Poly6_reg[6]  ( .D(n9687), .CP(clk), .CD(n18343), .Q(
        poly6_shifted[16]) );
  CFD2QXL \Poly6_reg[5]  ( .D(n9688), .CP(clk), .CD(n18344), .Q(
        poly6_shifted[15]) );
  CFD2QXL \Poly15_reg[34]  ( .D(n9603), .CP(clk), .CD(n18344), .Q(
        poly15_shifted[49]) );
  CFD2QXL \Poly15_reg[44]  ( .D(n9593), .CP(clk), .CD(n18345), .Q(
        poly15_shifted[59]) );
  CFD2QXL \Poly15_reg[39]  ( .D(n9598), .CP(clk), .CD(n18346), .Q(
        poly15_shifted[54]) );
  CFD2QXL \Poly1_reg[33]  ( .D(n9324), .CP(clk), .CD(n18358), .Q(
        poly1_shifted[44]) );
  CFD2QXL \Poly1_reg[66]  ( .D(n9291), .CP(clk), .CD(n18358), .Q(
        poly1_shifted[77]) );
  CFD2QXL \Poly1_reg[209]  ( .D(n9148), .CP(clk), .CD(n18359), .Q(
        poly1_shifted[220]) );
  CFD2QXL \Poly1_reg[242]  ( .D(n9115), .CP(clk), .CD(n18359), .Q(
        poly1_shifted[253]) );
  CFD2QXL \Poly1_reg[241]  ( .D(n9116), .CP(clk), .CD(n18360), .Q(
        poly1_shifted[252]) );
  CFD2QXL \Poly1_reg[240]  ( .D(n9117), .CP(clk), .CD(n18361), .Q(
        poly1_shifted[251]) );
  CFD2QXL \Poly1_reg[69]  ( .D(n9288), .CP(clk), .CD(n18362), .Q(
        poly1_shifted[80]) );
  CFD2QXL \Poly1_reg[35]  ( .D(n9322), .CP(clk), .CD(n18363), .Q(
        poly1_shifted[46]) );
  CFD2QXL \Poly1_reg[68]  ( .D(n9289), .CP(clk), .CD(n18363), .Q(
        poly1_shifted[79]) );
  CFD2QXL \Poly1_reg[167]  ( .D(n9190), .CP(clk), .CD(n18364), .Q(
        poly1_shifted[178]) );
  CFD2QXL \Poly1_reg[211]  ( .D(n9146), .CP(clk), .CD(n18364), .Q(
        poly1_shifted[222]) );
  CFD2QXL \Poly1_reg[238]  ( .D(n9119), .CP(clk), .CD(n18364), .Q(
        poly1_shifted[249]) );
  CFD2QXL \Poly1_reg[210]  ( .D(n9147), .CP(clk), .CD(n18254), .Q(
        poly1_shifted[221]) );
  CFD2QXL \Poly1_reg[237]  ( .D(n9120), .CP(clk), .CD(n18254), .Q(
        poly1_shifted[248]) );
  CFD2QXL \Poly1_reg[32]  ( .D(n9325), .CP(clk), .CD(n18366), .Q(
        poly1_shifted[43]) );
  CFD2QXL \Poly1_reg[65]  ( .D(n9292), .CP(clk), .CD(n18366), .Q(
        poly1_shifted[76]) );
  CFD2QXL \Poly1_reg[164]  ( .D(n9193), .CP(clk), .CD(n18367), .Q(
        poly1_shifted[175]) );
  CFD2QXL \Poly1_reg[246]  ( .D(n9111), .CP(clk), .CD(n18367), .Q(
        poly1_shifted[257]) );
  CFD2QXL \Poly1_reg[64]  ( .D(n9293), .CP(clk), .CD(n18368), .Q(
        poly1_shifted[75]) );
  CFD2QXL \Poly1_reg[218]  ( .D(n9139), .CP(clk), .CD(n18369), .Q(
        poly1_shifted[229]) );
  CFD2QXL \Poly1_reg[41]  ( .D(n9316), .CP(clk), .CD(n18370), .Q(
        poly1_shifted[52]) );
  CFD2QXL \Poly1_reg[74]  ( .D(n9283), .CP(clk), .CD(n18370), .Q(
        poly1_shifted[85]) );
  CFD2QXL \Poly1_reg[162]  ( .D(n9195), .CP(clk), .CD(n18370), .Q(
        poly1_shifted[173]) );
  CFD2QXL \Poly1_reg[217]  ( .D(n9140), .CP(clk), .CD(n18371), .Q(
        poly1_shifted[228]) );
  CFD2QXL \Poly1_reg[40]  ( .D(n9317), .CP(clk), .CD(n18372), .Q(
        poly1_shifted[51]) );
  CFD2QXL \Poly1_reg[172]  ( .D(n9185), .CP(clk), .CD(n18372), .Q(
        poly1_shifted[183]) );
  CFD2QXL \Poly1_reg[170]  ( .D(n9187), .CP(clk), .CD(n18373), .Q(
        poly1_shifted[181]) );
  CFD2QXL \Poly1_reg[214]  ( .D(n9143), .CP(clk), .CD(n18374), .Q(
        poly1_shifted[225]) );
  CFD2QXL \Poly1_reg[216]  ( .D(n9141), .CP(clk), .CD(n18374), .Q(
        poly1_shifted[227]) );
  CFD2QXL \Poly1_reg[243]  ( .D(n9114), .CP(clk), .CD(n18374), .Q(
        poly1_shifted[254]) );
  CFD2QXL \Poly1_reg[39]  ( .D(n9318), .CP(clk), .CD(n18374), .Q(
        poly1_shifted[50]) );
  CFD2QXL \Poly1_reg[72]  ( .D(n9285), .CP(clk), .CD(n18375), .Q(
        poly1_shifted[83]) );
  CFD2QXL \Poly1_reg[171]  ( .D(n9186), .CP(clk), .CD(n18375), .Q(
        poly1_shifted[182]) );
  CFD2QXL \Poly1_reg[37]  ( .D(n9320), .CP(clk), .CD(n18375), .Q(
        poly1_shifted[48]) );
  CFD2QXL \Poly1_reg[169]  ( .D(n9188), .CP(clk), .CD(n18376), .Q(
        poly1_shifted[180]) );
  CFD2QXL \Poly1_reg[213]  ( .D(n9144), .CP(clk), .CD(n18376), .Q(
        poly1_shifted[224]) );
  CFD2QXL \Poly1_reg[168]  ( .D(n9189), .CP(clk), .CD(n18377), .Q(
        poly1_shifted[179]) );
  CFD2QXL \Poly1_reg[215]  ( .D(n9142), .CP(clk), .CD(n18377), .Q(
        poly1_shifted[226]) );
  CFD2QXL \Poly3_reg[11]  ( .D(n8929), .CP(clk), .CD(n18384), .Q(
        poly3_shifted[25]) );
  CFD2QXL \Poly4_reg[15]  ( .D(n8841), .CP(clk), .CD(n18256), .Q(
        poly4_shifted[32]) );
  CFD2QXL \Poly4_reg[6]  ( .D(n8850), .CP(clk), .CD(n18256), .Q(
        poly4_shifted[23]) );
  CFD2QXL \Poly4_reg[5]  ( .D(n8851), .CP(clk), .CD(n18386), .Q(
        poly4_shifted[22]) );
  CFD2QXL \Poly4_reg[1]  ( .D(n8855), .CP(clk), .CD(n18386), .Q(
        poly4_shifted[18]) );
  CFD2QXL \Poly12_reg[98]  ( .D(n10434), .CP(clk), .CD(n18292), .Q(
        poly12_shifted[114]) );
  CFD2QXL \Poly12_reg[102]  ( .D(n10430), .CP(clk), .CD(n18293), .Q(
        poly12_shifted[118]) );
  CFD2QXL \Poly12_reg[104]  ( .D(n10428), .CP(clk), .CD(n18293), .Q(
        poly12_shifted[120]) );
  CFD2QXL \Poly12_reg[99]  ( .D(n10433), .CP(clk), .CD(n18294), .Q(
        poly12_shifted[115]) );
  CFD2QXL \Poly12_reg[101]  ( .D(n10431), .CP(clk), .CD(n18294), .Q(
        poly12_shifted[117]) );
  CFD2QXL \Poly12_reg[103]  ( .D(n10429), .CP(clk), .CD(n18295), .Q(
        poly12_shifted[119]) );
  CFD2QXL \Poly12_reg[107]  ( .D(n10425), .CP(clk), .CD(n18296), .Q(
        poly12_shifted[123]) );
  CFD2QXL \Poly12_reg[109]  ( .D(n10423), .CP(clk), .CD(n18297), .Q(
        poly12_shifted[125]) );
  CFD2QXL \Poly13_reg[482]  ( .D(n10578), .CP(clk), .CD(n18278), .Q(
        poly13_shifted[496]) );
  CFD2QXL \Poly13_reg[93]  ( .D(n10967), .CP(clk), .CD(n18281), .Q(
        poly13_shifted[107]) );
  CFD2QXL \Poly13_reg[33]  ( .D(n11027), .CP(clk), .CD(n18257), .Q(
        poly13_shifted[47]) );
  CFD2QXL \Poly14_reg[232]  ( .D(n10173), .CP(clk), .CD(n18303), .Q(
        poly14_shifted[248]) );
  CFD2QXL \Poly14_reg[149]  ( .D(n10256), .CP(clk), .CD(n18305), .Q(
        poly14_shifted[165]) );
  CFD2QXL \Poly6_reg[9]  ( .D(n9684), .CP(clk), .CD(n18342), .Q(
        poly6_shifted[19]) );
  CFD2QXL \Poly0_reg[36]  ( .D(n9541), .CP(clk), .CD(n18347), .Q(
        poly0_shifted[54]) );
  CFD2QXL \Poly0_reg[39]  ( .D(n9538), .CP(clk), .CD(n18349), .Q(
        poly0_shifted[57]) );
  CFD2QXL \Poly0_reg[129]  ( .D(n9448), .CP(clk), .CD(n18350), .Q(
        poly0_shifted[147]) );
  CFD2QXL \Poly0_reg[26]  ( .D(n9551), .CP(clk), .CD(n18350), .Q(
        poly0_shifted[44]) );
  CFD2QXL \Poly0_reg[23]  ( .D(n9554), .CP(clk), .CD(n18350), .Q(
        poly0_shifted[41]) );
  CFD2QXL \Poly0_reg[131]  ( .D(n9446), .CP(clk), .CD(n18351), .Q(
        poly0_shifted[149]) );
  CFD2QXL \Poly0_reg[30]  ( .D(n9547), .CP(clk), .CD(n18352), .Q(
        poly0_shifted[48]) );
  CFD2QXL \Poly0_reg[27]  ( .D(n9550), .CP(clk), .CD(n18352), .Q(
        poly0_shifted[45]) );
  CFD2QXL \Poly0_reg[32]  ( .D(n9545), .CP(clk), .CD(n18353), .Q(
        poly0_shifted[50]) );
  CFD2QXL \Poly0_reg[29]  ( .D(n9548), .CP(clk), .CD(n18353), .Q(
        poly0_shifted[47]) );
  CFD2QXL \Poly0_reg[137]  ( .D(n9440), .CP(clk), .CD(n18353), .Q(
        poly0_shifted[155]) );
  CFD2QXL \Poly0_reg[33]  ( .D(n9544), .CP(clk), .CD(n18355), .Q(
        poly0_shifted[51]) );
  CFD2QXL \Poly0_reg[38]  ( .D(n9539), .CP(clk), .CD(n18355), .Q(
        poly0_shifted[56]) );
  CFD2QXL \Poly0_reg[136]  ( .D(n9441), .CP(clk), .CD(n18356), .Q(
        poly0_shifted[154]) );
  CFD2QXL \Poly0_reg[35]  ( .D(n9542), .CP(clk), .CD(n18356), .Q(
        poly0_shifted[53]) );
  CFD2QXL \Poly0_reg[40]  ( .D(n9537), .CP(clk), .CD(n18356), .Q(
        poly0_shifted[58]) );
  CFD2QXL \Poly0_reg[130]  ( .D(n9447), .CP(clk), .CD(n18357), .Q(
        poly0_shifted[148]) );
  CFD2QXL \Poly0_reg[138]  ( .D(n9439), .CP(clk), .CD(n18357), .Q(
        poly0_shifted[156]) );
  CFD2QXL \Poly0_reg[24]  ( .D(n9553), .CP(clk), .CD(n18357), .Q(
        poly0_shifted[42]) );
  CFD2QXL \Poly3_reg[66]  ( .D(n8874), .CP(clk), .CD(n18382), .Q(
        poly3_shifted[80]) );
  CFD2QXL \Poly5_reg[14]  ( .D(n11512), .CP(clk), .CD(n18257), .Q(
        poly5_shifted[28]) );
  CFD2QXL \Poly5_reg[16]  ( .D(n11510), .CP(clk), .CD(n18258), .Q(
        poly5_shifted[30]) );
  CFD2QXL \Poly5_reg[13]  ( .D(n11513), .CP(clk), .CD(n18259), .Q(
        poly5_shifted[27]) );
  CFD2QXL \Poly5_reg[9]  ( .D(n11517), .CP(clk), .CD(n18257), .Q(
        poly5_shifted[23]) );
  CFD2QXL \Poly5_reg[15]  ( .D(n11511), .CP(clk), .CD(n18260), .Q(
        poly5_shifted[29]) );
  CFD2QXL \Poly13_reg[63]  ( .D(n10997), .CP(clk), .CD(n18285), .Q(
        poly13_shifted[77]) );
  CFD2QXL \Poly14_reg[31]  ( .D(n10374), .CP(clk), .CD(n18305), .Q(
        poly14_shifted[47]) );
  CFD2QXL \Poly0_reg[127]  ( .D(n9450), .CP(clk), .CD(n18357), .Q(
        poly0_shifted[145]) );
  CFD2QXL \Poly5_reg[34]  ( .D(n11492), .CP(clk), .CD(n18257), .Q(
        poly5_shifted[48]) );
  CFD2QXL \Poly5_reg[25]  ( .D(n11501), .CP(clk), .CD(n18257), .Q(
        poly5_shifted[39]) );
  CFD2QXL \Poly5_reg[57]  ( .D(n11469), .CP(clk), .CD(n18260), .Q(
        poly5_shifted[71]) );
  CFD2QXL \Poly8_reg[38]  ( .D(n11363), .CP(clk), .CD(n18257), .Q(
        poly8_shifted[52]) );
  CFD2QXL \Poly8_reg[50]  ( .D(n11351), .CP(clk), .CD(n18257), .Q(
        poly8_shifted[64]) );
  CFD2QXL \Poly8_reg[47]  ( .D(n11354), .CP(clk), .CD(n18257), .Q(
        poly8_shifted[61]) );
  CFD2QXL \Poly8_reg[34]  ( .D(n11367), .CP(clk), .CD(n18257), .Q(
        poly8_shifted[48]) );
  CFD2QXL \Poly13_reg[86]  ( .D(n10974), .CP(clk), .CD(n18257), .Q(
        poly13_shifted[100]) );
  CFD2QXL \Poly14_reg[264]  ( .D(n10141), .CP(clk), .CD(n18303), .Q(
        poly14_shifted[280]) );
  CFD2QXL \Poly14_reg[133]  ( .D(n10272), .CP(clk), .CD(n18305), .Q(
        poly14_shifted[149]) );
  CFD2QXL \Poly9_reg[35]  ( .D(n11270), .CP(clk), .CD(n18257), .Q(
        poly9_shifted[46]) );
  CFD2QXL \Poly13_reg[409]  ( .D(n10651), .CP(clk), .CD(n18284), .Q(
        poly13_shifted[423]) );
  CFD2QXL \Poly13_reg[289]  ( .D(n10771), .CP(clk), .CD(n18288), .Q(
        poly13_shifted[303]) );
  CFD2QXL \Poly1_reg[73]  ( .D(n9284), .CP(clk), .CD(n18372), .Q(
        poly1_shifted[84]) );
  CFD2QXL \Poly4_reg[41]  ( .D(n8815), .CP(clk), .CD(n18385), .Q(Poly4[41]) );
  CFD2QXL \Poly4_reg[40]  ( .D(n8816), .CP(clk), .CD(n18386), .Q(Poly4[40]) );
  CFD2QXL \Poly5_reg[98]  ( .D(n11428), .CP(clk), .CD(n18257), .Q(Poly5[98])
         );
  CFD2QXL \Poly5_reg[99]  ( .D(n11427), .CP(clk), .CD(n18258), .Q(Poly5[99])
         );
  CFD2QXL \Poly5_reg[94]  ( .D(n11432), .CP(clk), .CD(n18260), .Q(Poly5[94])
         );
  CFD2QXL \Poly5_reg[100]  ( .D(n11426), .CP(clk), .CD(n18257), .Q(Poly5[100])
         );
  CFD2QXL \Poly12_reg[34]  ( .D(n10498), .CP(clk), .CD(n18298), .Q(Poly12[34])
         );
  CFD2QXL \Poly12_reg[33]  ( .D(n10499), .CP(clk), .CD(n18298), .Q(Poly12[33])
         );
  CFD2QXL \Poly12_reg[81]  ( .D(n10451), .CP(clk), .CD(n18299), .Q(Poly12[81])
         );
  CFD2QXL \Poly14_reg[193]  ( .D(n10212), .CP(clk), .CD(n18308), .Q(
        Poly14[193]) );
  CFD2QXL \Poly14_reg[214]  ( .D(n10191), .CP(clk), .CD(n18309), .Q(
        Poly14[214]) );
  CFD2QXL \Poly14_reg[209]  ( .D(n10196), .CP(clk), .CD(n18310), .Q(
        Poly14[209]) );
  CFD2QXL \Poly7_reg[192]  ( .D(n9912), .CP(clk), .CD(n18317), .Q(Poly7[192])
         );
  CFD2QXL \Poly7_reg[191]  ( .D(n9913), .CP(clk), .CD(n18328), .Q(Poly7[191])
         );
  CFD2QXL \Poly7_reg[194]  ( .D(n9910), .CP(clk), .CD(n18329), .Q(Poly7[194])
         );
  CFD2QXL \Poly7_reg[193]  ( .D(n9911), .CP(clk), .CD(n18331), .Q(Poly7[193])
         );
  CFD2QXL \Poly7_reg[190]  ( .D(n9914), .CP(clk), .CD(n18341), .Q(Poly7[190])
         );
  CFD2QXL \Poly6_reg[38]  ( .D(n9655), .CP(clk), .CD(n18343), .Q(Poly6[38]) );
  CFD2QXL \Poly6_reg[31]  ( .D(n9662), .CP(clk), .CD(n18343), .Q(Poly6[31]) );
  CFD2QXL \Poly2_reg[39]  ( .D(n8971), .CP(clk), .CD(n18380), .Q(Poly2[39]) );
  CFD2QXL \Poly3_reg[56]  ( .D(n8884), .CP(clk), .CD(n18380), .Q(Poly3[56]) );
  CFD2QXL \dataselector_reg[41]  ( .D(n8754), .CP(clk), .CD(n18257), .Q(
        dataselector[41]) );
  CFD2QXL \dataselector_reg[20]  ( .D(n8775), .CP(clk), .CD(n18388), .Q(
        dataselector[20]) );
  CFD2QXL \Poly14_reg[175]  ( .D(n10230), .CP(clk), .CD(n18306), .Q(
        Poly14[175]) );
  CFD2QXL \Poly7_reg[180]  ( .D(n9924), .CP(clk), .CD(n18317), .Q(Poly7[180])
         );
  CFD2QXL \Poly0_reg[18]  ( .D(n9559), .CP(clk), .CD(n18347), .Q(Poly0[18]) );
  CFD2QXL \Poly0_reg[14]  ( .D(n9563), .CP(clk), .CD(n18347), .Q(Poly0[14]) );
  CFD2QXL \Poly0_reg[16]  ( .D(n9561), .CP(clk), .CD(n18347), .Q(Poly0[16]) );
  CFD2QXL \Poly0_reg[8]  ( .D(n9569), .CP(clk), .CD(n18348), .Q(Poly0[8]) );
  CFD2QXL \Poly0_reg[12]  ( .D(n9565), .CP(clk), .CD(n18349), .Q(Poly0[12]) );
  CFD2QXL \Poly0_reg[21]  ( .D(n9556), .CP(clk), .CD(n18349), .Q(Poly0[21]) );
  CFD2QXL \Poly0_reg[5]  ( .D(n9572), .CP(clk), .CD(n18350), .Q(Poly0[5]) );
  CFD2QXL \Poly0_reg[167]  ( .D(n9410), .CP(clk), .CD(n18351), .Q(Poly0[167])
         );
  CFD2QXL \Poly0_reg[7]  ( .D(n9570), .CP(clk), .CD(n18351), .Q(Poly0[7]) );
  CFD2QXL \Poly0_reg[153]  ( .D(n9424), .CP(clk), .CD(n18352), .Q(Poly0[153])
         );
  CFD2QXL \Poly0_reg[155]  ( .D(n9422), .CP(clk), .CD(n18353), .Q(Poly0[155])
         );
  CFD2QXL \Poly0_reg[160]  ( .D(n9417), .CP(clk), .CD(n18354), .Q(Poly0[160])
         );
  CFD2QXL \Poly0_reg[13]  ( .D(n9564), .CP(clk), .CD(n18354), .Q(Poly0[13]) );
  CFD2QXL \Poly0_reg[15]  ( .D(n9562), .CP(clk), .CD(n18355), .Q(Poly0[15]) );
  CFD2QXL \Poly0_reg[159]  ( .D(n9418), .CP(clk), .CD(n18355), .Q(Poly0[159])
         );
  CFD2QXL \Poly0_reg[154]  ( .D(n9423), .CP(clk), .CD(n18356), .Q(Poly0[154])
         );
  CFD2QXL \Poly0_reg[17]  ( .D(n9560), .CP(clk), .CD(n18356), .Q(Poly0[17]) );
  CFD2QXL \Poly0_reg[166]  ( .D(n9411), .CP(clk), .CD(n18357), .Q(Poly0[166])
         );
  CFD2QXL \Poly0_reg[158]  ( .D(n9419), .CP(clk), .CD(n18358), .Q(Poly0[158])
         );
  CFD2QXL \dataselector_reg[39]  ( .D(n8756), .CP(clk), .CD(n18257), .Q(
        dataselector[39]) );
  CFD2QXL \dataselector_reg[16]  ( .D(n8779), .CP(clk), .CD(n18387), .Q(
        dataselector[16]) );
  CFD2QXL \dataselector_reg[22]  ( .D(n8773), .CP(clk), .CD(n18387), .Q(
        dataselector[22]) );
  CFD2QXL \dataselector_reg[29]  ( .D(n8766), .CP(clk), .CD(n18387), .Q(
        dataselector[29]) );
  CFD2QXL \Poly6_reg[10]  ( .D(n9683), .CP(clk), .CD(n18341), .Q(Poly6[10]) );
  CFD2QXL \Poly4_reg[19]  ( .D(n8837), .CP(clk), .CD(n18385), .Q(Poly4[19]) );
  CFD2QXL \Poly6_reg[22]  ( .D(n9671), .CP(clk), .CD(n18396), .Q(Poly6[22]) );
  CFD2QXL \dataselector_reg[7]  ( .D(n8788), .CP(clk), .CD(n18388), .Q(
        dataselector[7]) );
  CFD2QXL \Poly13_reg[165]  ( .D(n10895), .CP(clk), .CD(n18278), .Q(
        Poly13[165]) );
  CFD2QXL \Poly14_reg[171]  ( .D(n10234), .CP(clk), .CD(n18304), .Q(
        Poly14[171]) );
  CFD2QXL \Poly2_reg[48]  ( .D(n8962), .CP(clk), .CD(n18377), .Q(Poly2[48]) );
  CFD2QXL \Poly2_reg[32]  ( .D(n8978), .CP(clk), .CD(n18391), .Q(Poly2[32]) );
  CFD2QXL \Poly10_reg[17]  ( .D(n11086), .CP(clk), .CD(n18263), .Q(Poly10[17])
         );
  CFD2QXL \Poly0_reg[108]  ( .D(n9469), .CP(clk), .CD(n18347), .Q(Poly0[108])
         );
  CFD2QXL \Poly0_reg[117]  ( .D(n9460), .CP(clk), .CD(n18352), .Q(Poly0[117])
         );
  CFD2QXL \Poly0_reg[104]  ( .D(n9473), .CP(clk), .CD(n18353), .Q(Poly0[104])
         );
  CFD2QXL \Poly8_reg[9]  ( .D(n11392), .CP(clk), .CD(n18261), .Q(Poly8[9]) );
  CFD2QXL \Poly11_reg[29]  ( .D(n11160), .CP(clk), .CD(n18257), .Q(Poly11[29])
         );
  CFD2QXL \Poly8_reg[18]  ( .D(n11383), .CP(clk), .CD(n18257), .Q(
        poly8_shifted[32]) );
  CFD2QXL \Poly1_reg[36]  ( .D(n9321), .CP(clk), .CD(n18361), .Q(
        poly1_shifted[47]) );
  CFD2QXL \Poly6_reg[3]  ( .D(n9690), .CP(clk), .CD(n18343), .Q(Poly6[3]) );
  CFD2QXL \Poly11_reg[69]  ( .D(n11120), .CP(clk), .CD(n18257), .Q(Poly11[69])
         );
  CFD2QXL \Poly12_reg[57]  ( .D(n10475), .CP(clk), .CD(n18296), .Q(Poly12[57])
         );
  CFD2QXL \Poly2_reg[47]  ( .D(n8963), .CP(clk), .CD(n18390), .Q(Poly2[47]) );
  CFD2QXL \Poly12_reg[108]  ( .D(n10424), .CP(clk), .CD(n18294), .Q(
        poly12_shifted[124]) );
  CFD2QXL \Poly0_reg[146]  ( .D(n9431), .CP(clk), .CD(n18355), .Q(
        poly0_shifted[164]) );
  CFD2QXL \Poly5_reg[49]  ( .D(n11477), .CP(clk), .CD(n18259), .Q(
        poly5_shifted[63]) );
  CFD2QXL \Poly11_reg[77]  ( .D(n11112), .CP(clk), .CD(n18262), .Q(Poly11[77])
         );
  CFD2QXL \Poly15_reg[26]  ( .D(n9611), .CP(clk), .CD(n18346), .Q(Poly15[26])
         );
  CFD2QXL \Poly8_reg[14]  ( .D(n11387), .CP(clk), .CD(n18257), .Q(Poly8[14])
         );
  CFD2QXL \Poly8_reg[70]  ( .D(n11331), .CP(clk), .CD(n18257), .Q(Poly8[70])
         );
  CFD2QXL \Poly8_reg[72]  ( .D(n11329), .CP(clk), .CD(n18257), .Q(Poly8[72])
         );
  CFD2QXL \Poly8_reg[12]  ( .D(n11389), .CP(clk), .CD(n18257), .Q(Poly8[12])
         );
  CFD2QXL \Poly8_reg[71]  ( .D(n11330), .CP(clk), .CD(n18257), .Q(Poly8[71])
         );
  CFD2QXL \Poly8_reg[69]  ( .D(n11332), .CP(clk), .CD(n18261), .Q(Poly8[69])
         );
  CFD2QXL \Poly8_reg[80]  ( .D(n11321), .CP(clk), .CD(n18257), .Q(Poly8[80])
         );
  CFD2QXL \Poly8_reg[79]  ( .D(n11322), .CP(clk), .CD(n18257), .Q(Poly8[79])
         );
  CFD2QXL \Poly8_reg[4]  ( .D(n11397), .CP(clk), .CD(n18257), .Q(Poly8[4]) );
  CFD2QXL \Poly8_reg[77]  ( .D(n11324), .CP(clk), .CD(n18257), .Q(Poly8[77])
         );
  CFD2QXL \Poly9_reg[20]  ( .D(n11285), .CP(clk), .CD(n18257), .Q(Poly9[20])
         );
  CFD2QXL \Poly9_reg[21]  ( .D(n11284), .CP(clk), .CD(n18257), .Q(Poly9[21])
         );
  CFD2QXL \Poly9_reg[13]  ( .D(n11292), .CP(clk), .CD(n18257), .Q(Poly9[13])
         );
  CFD2QXL \Poly9_reg[90]  ( .D(n11215), .CP(clk), .CD(n18257), .Q(Poly9[90])
         );
  CFD2QXL \Poly9_reg[92]  ( .D(n11213), .CP(clk), .CD(n18257), .Q(Poly9[92])
         );
  CFD2QXL \Poly11_reg[30]  ( .D(n11159), .CP(clk), .CD(n18257), .Q(Poly11[30])
         );
  CFD2QXL \Poly11_reg[19]  ( .D(n11170), .CP(clk), .CD(n18257), .Q(Poly11[19])
         );
  CFD2QXL \Poly11_reg[26]  ( .D(n11163), .CP(clk), .CD(n18257), .Q(Poly11[26])
         );
  CFD2QXL \Poly11_reg[18]  ( .D(n11171), .CP(clk), .CD(n18257), .Q(Poly11[18])
         );
  CFD2QXL \Poly11_reg[31]  ( .D(n11158), .CP(clk), .CD(n18257), .Q(Poly11[31])
         );
  CFD2QXL \Poly11_reg[22]  ( .D(n11167), .CP(clk), .CD(n18257), .Q(Poly11[22])
         );
  CFD2QXL \Poly11_reg[62]  ( .D(n11127), .CP(clk), .CD(n18257), .Q(Poly11[62])
         );
  CFD2QXL \Poly11_reg[20]  ( .D(n11169), .CP(clk), .CD(n18257), .Q(Poly11[20])
         );
  CFD2QXL \Poly11_reg[37]  ( .D(n11152), .CP(clk), .CD(n18257), .Q(Poly11[37])
         );
  CFD2QXL \Poly11_reg[70]  ( .D(n11119), .CP(clk), .CD(n18257), .Q(Poly11[70])
         );
  CFD2QXL \Poly11_reg[27]  ( .D(n11162), .CP(clk), .CD(n18257), .Q(Poly11[27])
         );
  CFD2QXL \Poly11_reg[59]  ( .D(n11130), .CP(clk), .CD(n18262), .Q(Poly11[59])
         );
  CFD2QXL \Poly13_reg[280]  ( .D(n10780), .CP(clk), .CD(n18265), .Q(
        Poly13[280]) );
  CFD2QXL \Poly13_reg[156]  ( .D(n10904), .CP(clk), .CD(n18257), .Q(
        Poly13[156]) );
  CFD2QXL \Poly13_reg[269]  ( .D(n10791), .CP(clk), .CD(n18257), .Q(
        Poly13[269]) );
  CFD2QXL \Poly13_reg[167]  ( .D(n10893), .CP(clk), .CD(n18275), .Q(
        Poly13[167]) );
  CFD2QXL \Poly13_reg[166]  ( .D(n10894), .CP(clk), .CD(n18276), .Q(
        Poly13[166]) );
  CFD2QXL \Poly13_reg[279]  ( .D(n10781), .CP(clk), .CD(n18255), .Q(
        Poly13[279]) );
  CFD2QXL \Poly13_reg[278]  ( .D(n10782), .CP(clk), .CD(n18278), .Q(
        Poly13[278]) );
  CFD2QXL \Poly13_reg[391]  ( .D(n10669), .CP(clk), .CD(n18280), .Q(
        Poly13[391]) );
  CFD2QXL \Poly13_reg[390]  ( .D(n10670), .CP(clk), .CD(n18283), .Q(
        Poly13[390]) );
  CFD2QXL \Poly13_reg[389]  ( .D(n10671), .CP(clk), .CD(n18284), .Q(
        Poly13[389]) );
  CFD2QXL \Poly13_reg[160]  ( .D(n10900), .CP(clk), .CD(n18287), .Q(
        Poly13[160]) );
  CFD2QXL \Poly13_reg[399]  ( .D(n10661), .CP(clk), .CD(n18288), .Q(
        Poly13[399]) );
  CFD2QXL \Poly13_reg[159]  ( .D(n10901), .CP(clk), .CD(n18257), .Q(
        Poly13[159]) );
  CFD2QXL \Poly13_reg[271]  ( .D(n10789), .CP(clk), .CD(n18290), .Q(
        Poly13[271]) );
  CFD2QXL \Poly13_reg[397]  ( .D(n10663), .CP(clk), .CD(n18290), .Q(
        Poly13[397]) );
  CFD2QXL \Poly13_reg[272]  ( .D(n10788), .CP(clk), .CD(n18291), .Q(
        Poly13[272]) );
  CFD2QXL \Poly13_reg[400]  ( .D(n10660), .CP(clk), .CD(n18292), .Q(
        Poly13[400]) );
  CFD2QXL \Poly12_reg[21]  ( .D(n10511), .CP(clk), .CD(n18293), .Q(Poly12[21])
         );
  CFD2QXL \Poly12_reg[23]  ( .D(n10509), .CP(clk), .CD(n18293), .Q(Poly12[23])
         );
  CFD2QXL \Poly12_reg[20]  ( .D(n10512), .CP(clk), .CD(n18294), .Q(Poly12[20])
         );
  CFD2QXL \Poly12_reg[36]  ( .D(n10496), .CP(clk), .CD(n18294), .Q(Poly12[36])
         );
  CFD2QXL \Poly12_reg[22]  ( .D(n10510), .CP(clk), .CD(n18295), .Q(Poly12[22])
         );
  CFD2QXL \Poly12_reg[37]  ( .D(n10495), .CP(clk), .CD(n18295), .Q(Poly12[37])
         );
  CFD2QXL \Poly12_reg[53]  ( .D(n10479), .CP(clk), .CD(n18295), .Q(Poly12[53])
         );
  CFD2QXL \Poly12_reg[26]  ( .D(n10506), .CP(clk), .CD(n18295), .Q(Poly12[26])
         );
  CFD2QXL \Poly12_reg[60]  ( .D(n10472), .CP(clk), .CD(n18296), .Q(Poly12[60])
         );
  CFD2QXL \Poly12_reg[59]  ( .D(n10473), .CP(clk), .CD(n18296), .Q(Poly12[59])
         );
  CFD2QXL \Poly12_reg[30]  ( .D(n10502), .CP(clk), .CD(n18297), .Q(Poly12[30])
         );
  CFD2QXL \Poly12_reg[61]  ( .D(n10471), .CP(clk), .CD(n18297), .Q(Poly12[61])
         );
  CFD2QXL \Poly12_reg[63]  ( .D(n10469), .CP(clk), .CD(n18298), .Q(Poly12[63])
         );
  CFD2QXL \Poly12_reg[84]  ( .D(n10448), .CP(clk), .CD(n18298), .Q(Poly12[84])
         );
  CFD2QXL \Poly12_reg[65]  ( .D(n10467), .CP(clk), .CD(n18299), .Q(Poly12[65])
         );
  CFD2QXL \Poly12_reg[56]  ( .D(n10476), .CP(clk), .CD(n18299), .Q(Poly12[56])
         );
  CFD2QXL \Poly14_reg[173]  ( .D(n10232), .CP(clk), .CD(n18301), .Q(
        Poly14[173]) );
  CFD2QXL \Poly14_reg[165]  ( .D(n10240), .CP(clk), .CD(n18305), .Q(
        Poly14[165]) );
  CFD2QXL \Poly14_reg[201]  ( .D(n10204), .CP(clk), .CD(n18307), .Q(
        Poly14[201]) );
  CFD2QXL \Poly14_reg[204]  ( .D(n10201), .CP(clk), .CD(n18308), .Q(
        Poly14[204]) );
  CFD2QXL \Poly14_reg[197]  ( .D(n10208), .CP(clk), .CD(n18310), .Q(
        Poly14[197]) );
  CFD2QXL \Poly14_reg[207]  ( .D(n10198), .CP(clk), .CD(n18311), .Q(
        Poly14[207]) );
  CFD2QXL \Poly14_reg[180]  ( .D(n10225), .CP(clk), .CD(n18312), .Q(
        Poly14[180]) );
  CFD2QXL \Poly14_reg[196]  ( .D(n10209), .CP(clk), .CD(n18312), .Q(
        Poly14[196]) );
  CFD2QXL \Poly14_reg[212]  ( .D(n10193), .CP(clk), .CD(n18312), .Q(
        Poly14[212]) );
  CFD2QXL \Poly14_reg[174]  ( .D(n10231), .CP(clk), .CD(n18313), .Q(
        Poly14[174]) );
  CFD2QXL \Poly14_reg[168]  ( .D(n10237), .CP(clk), .CD(n18315), .Q(
        Poly14[168]) );
  CFD2QXL \Poly14_reg[206]  ( .D(n10199), .CP(clk), .CD(n18316), .Q(
        Poly14[206]) );
  CFD2QXL \Poly7_reg[19]  ( .D(n10085), .CP(clk), .CD(n18323), .Q(Poly7[19])
         );
  CFD2QXL \Poly7_reg[233]  ( .D(n9871), .CP(clk), .CD(n18324), .Q(Poly7[233])
         );
  CFD2QXL \Poly7_reg[189]  ( .D(n9915), .CP(clk), .CD(n18326), .Q(Poly7[189])
         );
  CFD2QXL \Poly7_reg[184]  ( .D(n9920), .CP(clk), .CD(n18329), .Q(Poly7[184])
         );
  CFD2QXL \Poly7_reg[49]  ( .D(n10055), .CP(clk), .CD(n18331), .Q(Poly7[49])
         );
  CFD2QXL \Poly7_reg[183]  ( .D(n9921), .CP(clk), .CD(n18335), .Q(Poly7[183])
         );
  CFD2QXL \Poly7_reg[188]  ( .D(n9916), .CP(clk), .CD(n18335), .Q(Poly7[188])
         );
  CFD2QXL \Poly7_reg[239]  ( .D(n9865), .CP(clk), .CD(n18336), .Q(Poly7[239])
         );
  CFD2QXL \Poly7_reg[241]  ( .D(n9863), .CP(clk), .CD(n18339), .Q(Poly7[241])
         );
  CFD2QXL \Poly0_reg[152]  ( .D(n9425), .CP(clk), .CD(n18354), .Q(Poly0[152])
         );
  CFD2QXL \Poly1_reg[208]  ( .D(n9149), .CP(clk), .CD(n18367), .Q(Poly1[208])
         );
  CFD2QXL \Poly2_reg[19]  ( .D(n8991), .CP(clk), .CD(n18378), .Q(Poly2[19]) );
  CFD2QXL \Poly2_reg[18]  ( .D(n8992), .CP(clk), .CD(n18378), .Q(Poly2[18]) );
  CFD2QXL \Poly2_reg[20]  ( .D(n8990), .CP(clk), .CD(n18378), .Q(Poly2[20]) );
  CFD2QXL \Poly2_reg[27]  ( .D(n8983), .CP(clk), .CD(n18379), .Q(Poly2[27]) );
  CFD2QXL \Poly3_reg[40]  ( .D(n8900), .CP(clk), .CD(n18381), .Q(Poly3[40]) );
  CFD2QXL \Poly3_reg[43]  ( .D(n8897), .CP(clk), .CD(n18382), .Q(Poly3[43]) );
  CFD2QXL \Poly3_reg[38]  ( .D(n8902), .CP(clk), .CD(n18383), .Q(Poly3[38]) );
  CFD2QXL \Poly4_reg[18]  ( .D(n8838), .CP(clk), .CD(n18386), .Q(Poly4[18]) );
  CFD2QXL \Poly0_reg[173]  ( .D(n9404), .CP(clk), .CD(n18351), .Q(
        poly0_shifted[191]) );
  CFD2QXL \Poly5_reg[72]  ( .D(n11454), .CP(clk), .CD(n18258), .Q(
        poly5_shifted[86]) );
  CFD2QXL \Poly5_reg[78]  ( .D(n11448), .CP(clk), .CD(n18257), .Q(Poly5[78])
         );
  CFD2QXL \Poly5_reg[69]  ( .D(n11457), .CP(clk), .CD(n18259), .Q(
        poly5_shifted[83]) );
  CFD2QXL \Poly5_reg[48]  ( .D(n11478), .CP(clk), .CD(n18257), .Q(
        poly5_shifted[62]) );
  CFD2QXL \Poly5_reg[67]  ( .D(n11459), .CP(clk), .CD(n18257), .Q(
        poly5_shifted[81]) );
  CFD2QXL \Poly5_reg[54]  ( .D(n11472), .CP(clk), .CD(n18257), .Q(
        poly5_shifted[68]) );
  CFD2QXL \Poly5_reg[46]  ( .D(n11480), .CP(clk), .CD(n18257), .Q(
        poly5_shifted[60]) );
  CFD2QXL \Poly5_reg[65]  ( .D(n11461), .CP(clk), .CD(n18260), .Q(
        poly5_shifted[79]) );
  CFD2QXL \Poly5_reg[71]  ( .D(n11455), .CP(clk), .CD(n18257), .Q(
        poly5_shifted[85]) );
  CFD2QXL \Poly15_reg[42]  ( .D(n9595), .CP(clk), .CD(n18345), .Q(
        poly15_shifted[57]) );
  CFD2QXL \Poly15_reg[43]  ( .D(n9594), .CP(clk), .CD(n18396), .Q(
        poly15_shifted[58]) );
  CFD2QXL \Poly15_reg[36]  ( .D(n9601), .CP(clk), .CD(n18256), .Q(
        poly15_shifted[51]) );
  CFD2QXL \Poly0_reg[98]  ( .D(n9479), .CP(clk), .CD(n18350), .Q(
        poly0_shifted[116]) );
  CFD2QXL \Poly0_reg[97]  ( .D(n9480), .CP(clk), .CD(n18352), .Q(
        poly0_shifted[115]) );
  CFD2QXL \Poly0_reg[102]  ( .D(n9475), .CP(clk), .CD(n18352), .Q(
        poly0_shifted[120]) );
  CFD2QXL \Poly0_reg[99]  ( .D(n9478), .CP(clk), .CD(n18352), .Q(
        poly0_shifted[117]) );
  CFD2QXL \dataselector_reg[35]  ( .D(n8760), .CP(clk), .CD(n18388), .Q(
        dataselector[35]) );
  CFD2QXL \dataselector_reg[45]  ( .D(n8750), .CP(clk), .CD(n18387), .Q(
        dataselector[45]) );
  CFD2QXL \dataselector_reg[43]  ( .D(n8752), .CP(clk), .CD(n18387), .Q(
        dataselector[43]) );
  CFD2QXL \Poly0_reg[145]  ( .D(n9432), .CP(clk), .CD(n18394), .Q(
        poly0_shifted[163]) );
  CFD2QXL \Poly6_reg[39]  ( .D(n9654), .CP(clk), .CD(n18342), .Q(Poly6[39]) );
  CFD2QXL \Poly10_reg[11]  ( .D(n11092), .CP(clk), .CD(n18400), .Q(Poly10[11])
         );
  CFD2QXL \Poly0_reg[139]  ( .D(n9438), .CP(clk), .CD(n18354), .Q(
        poly0_shifted[157]) );
  CFD2QXL \Poly5_reg[47]  ( .D(n11479), .CP(clk), .CD(n18257), .Q(
        poly5_shifted[61]) );
  CFD2QXL \Poly5_reg[75]  ( .D(n11451), .CP(clk), .CD(n18257), .Q(
        poly5_shifted[89]) );
  CFD2QXL \Poly5_reg[39]  ( .D(n11487), .CP(clk), .CD(n18257), .Q(
        poly5_shifted[53]) );
  CFD2QXL \Poly5_reg[37]  ( .D(n11489), .CP(clk), .CD(n18260), .Q(
        poly5_shifted[51]) );
  CFD2QXL \Poly11_reg[64]  ( .D(n11125), .CP(clk), .CD(n18257), .Q(Poly11[64])
         );
  CFD2QXL \Poly15_reg[49]  ( .D(n9588), .CP(clk), .CD(n18344), .Q(Poly15[49])
         );
  CFD2QXL \Poly15_reg[48]  ( .D(n9589), .CP(clk), .CD(n18346), .Q(Poly15[48])
         );
  CFD2QXL \Poly15_reg[58]  ( .D(n9579), .CP(clk), .CD(n18256), .Q(Poly15[58])
         );
  CFD2QXL \Poly3_reg[82]  ( .D(n8858), .CP(clk), .CD(n18381), .Q(Poly3[82]) );
  CFD2QXL \Poly3_reg[71]  ( .D(n8869), .CP(clk), .CD(n18382), .Q(Poly3[71]) );
  CFD2QXL \Poly4_reg[29]  ( .D(n8827), .CP(clk), .CD(n18385), .Q(Poly4[29]) );
  CFD2QXL \Poly15_reg[23]  ( .D(n9614), .CP(clk), .CD(n18345), .Q(Poly15[23])
         );
  CFD2QXL \Poly2_reg[22]  ( .D(n8988), .CP(clk), .CD(n18379), .Q(Poly2[22]) );
  CFD2QXL \Poly4_reg[31]  ( .D(n8825), .CP(clk), .CD(n18386), .Q(Poly4[31]) );
  CFD2QXL \Poly8_reg[15]  ( .D(n11386), .CP(clk), .CD(n18257), .Q(Poly8[15])
         );
  CFD2QXL \Poly8_reg[13]  ( .D(n11388), .CP(clk), .CD(n18257), .Q(Poly8[13])
         );
  CFD2QXL \Poly8_reg[11]  ( .D(n11390), .CP(clk), .CD(n18257), .Q(Poly8[11])
         );
  CFD2QXL \Poly8_reg[10]  ( .D(n11391), .CP(clk), .CD(n18257), .Q(Poly8[10])
         );
  CFD2QXL \Poly8_reg[7]  ( .D(n11394), .CP(clk), .CD(n18257), .Q(Poly8[7]) );
  CFD2QXL \Poly8_reg[6]  ( .D(n11395), .CP(clk), .CD(n18257), .Q(Poly8[6]) );
  CFD2QXL \Poly8_reg[5]  ( .D(n11396), .CP(clk), .CD(n18257), .Q(Poly8[5]) );
  CFD2QXL \Poly9_reg[16]  ( .D(n11289), .CP(clk), .CD(n18257), .Q(Poly9[16])
         );
  CFD2QXL \Poly9_reg[18]  ( .D(n11287), .CP(clk), .CD(n18257), .Q(Poly9[18])
         );
  CFD2QXL \Poly9_reg[19]  ( .D(n11286), .CP(clk), .CD(n18257), .Q(Poly9[19])
         );
  CFD2QXL \Poly11_reg[41]  ( .D(n11148), .CP(clk), .CD(n18257), .Q(Poly11[41])
         );
  CFD2QXL \Poly11_reg[47]  ( .D(n11142), .CP(clk), .CD(n18257), .Q(Poly11[47])
         );
  CFD2QXL \Poly11_reg[44]  ( .D(n11145), .CP(clk), .CD(n18262), .Q(Poly11[44])
         );
  CFD2QXL \Poly12_reg[25]  ( .D(n10507), .CP(clk), .CD(n18293), .Q(Poly12[25])
         );
  CFD2QXL \Poly12_reg[24]  ( .D(n10508), .CP(clk), .CD(n18295), .Q(Poly12[24])
         );
  CFD2QXL \Poly12_reg[55]  ( .D(n10477), .CP(clk), .CD(n18295), .Q(Poly12[55])
         );
  CFD2QXL \Poly12_reg[62]  ( .D(n10470), .CP(clk), .CD(n18297), .Q(Poly12[62])
         );
  CFD2QXL \Poly12_reg[52]  ( .D(n10480), .CP(clk), .CD(n18297), .Q(Poly12[52])
         );
  CFD2QXL \Poly12_reg[66]  ( .D(n10466), .CP(clk), .CD(n18298), .Q(Poly12[66])
         );
  CFD2QXL \Poly14_reg[208]  ( .D(n10197), .CP(clk), .CD(n18254), .Q(
        Poly14[208]) );
  CFD2QXL \Poly14_reg[203]  ( .D(n10202), .CP(clk), .CD(n18309), .Q(
        Poly14[203]) );
  CFD2QXL \Poly14_reg[202]  ( .D(n10203), .CP(clk), .CD(n18311), .Q(
        Poly14[202]) );
  CFD2QXL \Poly14_reg[200]  ( .D(n10205), .CP(clk), .CD(n18315), .Q(
        Poly14[200]) );
  CFD2QXL \Poly14_reg[199]  ( .D(n10206), .CP(clk), .CD(n18316), .Q(
        Poly14[199]) );
  CFD2QXL \Poly7_reg[186]  ( .D(n9918), .CP(clk), .CD(n18332), .Q(Poly7[186])
         );
  CFD2QXL \Poly7_reg[185]  ( .D(n9919), .CP(clk), .CD(n18338), .Q(Poly7[185])
         );
  CFD2QXL \Poly15_reg[19]  ( .D(n9618), .CP(clk), .CD(n18345), .Q(Poly15[19])
         );
  CFD2QXL \Poly15_reg[18]  ( .D(n9619), .CP(clk), .CD(n18346), .Q(Poly15[18])
         );
  CFD2QXL \Poly15_reg[20]  ( .D(n9617), .CP(clk), .CD(n18346), .Q(Poly15[20])
         );
  CFD2QXL \Poly2_reg[23]  ( .D(n8987), .CP(clk), .CD(n18378), .Q(Poly2[23]) );
  CFD2QXL \Poly3_reg[37]  ( .D(n8903), .CP(clk), .CD(n18381), .Q(Poly3[37]) );
  CFD2QXL \Poly3_reg[44]  ( .D(n8896), .CP(clk), .CD(n18383), .Q(Poly3[44]) );
  CFD2QXL \Poly0_reg[46]  ( .D(n9531), .CP(clk), .CD(n18395), .Q(
        poly0_shifted[64]) );
  CFD2QXL \Poly5_reg[104]  ( .D(n11422), .CP(clk), .CD(n18257), .Q(
        poly5_shifted[118]) );
  CFD2QXL \Poly8_reg[57]  ( .D(n11344), .CP(clk), .CD(n18257), .Q(
        poly8_shifted[71]) );
  CFD2QXL \Poly8_reg[51]  ( .D(n11350), .CP(clk), .CD(n18257), .Q(
        poly8_shifted[65]) );
  CFD2QXL \Poly9_reg[28]  ( .D(n11277), .CP(clk), .CD(n18257), .Q(
        poly9_shifted[39]) );
  CFD2QXL \Poly11_reg[6]  ( .D(n11183), .CP(clk), .CD(n18257), .Q(
        poly11_shifted[21]) );
  CFD2QXL \Poly11_reg[12]  ( .D(n11177), .CP(clk), .CD(n18257), .Q(
        poly11_shifted[27]) );
  CFD2QXL \Poly13_reg[28]  ( .D(n11032), .CP(clk), .CD(n18264), .Q(
        poly13_shifted[42]) );
  CFD2QXL \Poly13_reg[32]  ( .D(n11028), .CP(clk), .CD(n18266), .Q(
        poly13_shifted[46]) );
  CFD2QXL \Poly13_reg[16]  ( .D(n11044), .CP(clk), .CD(n18269), .Q(
        poly13_shifted[30]) );
  CFD2QXL \Poly13_reg[1]  ( .D(n11059), .CP(clk), .CD(n18270), .Q(
        poly13_shifted[15]) );
  CFD2QXL \Poly13_reg[43]  ( .D(n11017), .CP(clk), .CD(n18270), .Q(
        poly13_shifted[57]) );
  CFD2QXL \Poly13_reg[13]  ( .D(n11047), .CP(clk), .CD(n18274), .Q(
        poly13_shifted[27]) );
  CFD2QXL \Poly13_reg[41]  ( .D(n11019), .CP(clk), .CD(n18274), .Q(
        poly13_shifted[55]) );
  CFD2QXL \Poly13_reg[25]  ( .D(n11035), .CP(clk), .CD(n18277), .Q(
        poly13_shifted[39]) );
  CFD2QXL \Poly12_reg[71]  ( .D(n10461), .CP(clk), .CD(n18295), .Q(
        poly12_shifted[87]) );
  CFD2QXL \Poly14_reg[224]  ( .D(n10181), .CP(clk), .CD(n18254), .Q(
        poly14_shifted[240]) );
  CFD2QXL \Poly14_reg[39]  ( .D(n10366), .CP(clk), .CD(n18302), .Q(
        poly14_shifted[55]) );
  CFD2QXL \Poly14_reg[215]  ( .D(n10190), .CP(clk), .CD(n18310), .Q(
        poly14_shifted[231]) );
  CFD2QXL \Poly7_reg[197]  ( .D(n9907), .CP(clk), .CD(n18324), .Q(
        poly7_shifted[209]) );
  CFD2QXL \Poly7_reg[104]  ( .D(n10000), .CP(clk), .CD(n18335), .Q(
        poly7_shifted[116]) );
  CFD2QXL \Poly7_reg[198]  ( .D(n9906), .CP(clk), .CD(n18335), .Q(
        poly7_shifted[210]) );
  CFD2QXL \Poly7_reg[327]  ( .D(n9777), .CP(clk), .CD(n18339), .Q(
        poly7_shifted[339]) );
  CFD2QXL \Poly7_reg[351]  ( .D(n9753), .CP(clk), .CD(n18339), .Q(
        poly7_shifted[363]) );
  CFD2QXL \Poly7_reg[115]  ( .D(n9989), .CP(clk), .CD(n18340), .Q(
        poly7_shifted[127]) );
  CFD2QXL \Poly7_reg[199]  ( .D(n9905), .CP(clk), .CD(n18340), .Q(
        poly7_shifted[211]) );
  CFD2QXL \Poly1_reg[47]  ( .D(n9310), .CP(clk), .CD(n18361), .Q(
        poly1_shifted[58]) );
  CFD2QXL \Poly1_reg[290]  ( .D(n9067), .CP(clk), .CD(n18367), .Q(
        poly1_shifted[301]) );
  CFD2QXL \Poly1_reg[42]  ( .D(n9315), .CP(clk), .CD(n18368), .Q(
        poly1_shifted[53]) );
  CFD2QXL \Poly1_reg[267]  ( .D(n9090), .CP(clk), .CD(n18369), .Q(
        poly1_shifted[278]) );
  CFD2QXL \Poly1_reg[49]  ( .D(n9308), .CP(clk), .CD(n18373), .Q(
        poly1_shifted[60]) );
  CFD2QXL \Poly4_reg[7]  ( .D(n8849), .CP(clk), .CD(n18385), .Q(
        poly4_shifted[24]) );
  CFD2QXL \Poly4_reg[10]  ( .D(n8846), .CP(clk), .CD(n18386), .Q(
        poly4_shifted[27]) );
  CFD2QXL \Poly6_reg[2]  ( .D(n9691), .CP(clk), .CD(n18342), .Q(Poly6[2]) );
  CFD2QXL \Poly3_reg[64]  ( .D(n8876), .CP(clk), .CD(n18384), .Q(
        poly3_shifted[78]) );
  CFD2QXL \Poly5_reg[0]  ( .D(n11526), .CP(clk), .CD(n18257), .Q(Poly5[0]) );
  CFD2QXL \Poly5_reg[3]  ( .D(n11523), .CP(clk), .CD(n18258), .Q(Poly5[3]) );
  CFD2QXL \Poly5_reg[4]  ( .D(n11522), .CP(clk), .CD(n18257), .Q(Poly5[4]) );
  CFD2QXL \dataselector_reg[17]  ( .D(n8778), .CP(clk), .CD(n18388), .Q(
        dataselector[17]) );
  CFD2QXL \dataselector_reg[9]  ( .D(n8786), .CP(clk), .CD(n18388), .Q(
        dataselector[9]) );
  CFD2QXL \scrambler_reg[8]  ( .D(n8708), .CP(clk), .CD(n18401), .Q(
        scrambler[8]) );
  CFD2QXL \Poly5_reg[83]  ( .D(n11443), .CP(clk), .CD(n18257), .Q(Poly5[83])
         );
  CFD2QXL \Poly5_reg[76]  ( .D(n11450), .CP(clk), .CD(n18257), .Q(Poly5[76])
         );
  CFD2QXL \Poly5_reg[81]  ( .D(n11445), .CP(clk), .CD(n18257), .Q(Poly5[81])
         );
  CFD2QXL \Poly5_reg[87]  ( .D(n11439), .CP(clk), .CD(n18257), .Q(Poly5[87])
         );
  CFD2QXL \Poly5_reg[88]  ( .D(n11438), .CP(clk), .CD(n18257), .Q(Poly5[88])
         );
  CFD2QXL \Poly5_reg[93]  ( .D(n11433), .CP(clk), .CD(n18260), .Q(Poly5[93])
         );
  CFD2QXL \Poly9_reg[14]  ( .D(n11291), .CP(clk), .CD(n18257), .Q(Poly9[14])
         );
  CFD2QXL \Poly14_reg[169]  ( .D(n10236), .CP(clk), .CD(n18307), .Q(
        Poly14[169]) );
  CFD2QXL \Poly14_reg[178]  ( .D(n10227), .CP(clk), .CD(n18316), .Q(
        Poly14[178]) );
  CFD2QXL \Poly7_reg[52]  ( .D(n10052), .CP(clk), .CD(n18328), .Q(Poly7[52])
         );
  CFD2QXL \Poly7_reg[58]  ( .D(n10046), .CP(clk), .CD(n18337), .Q(Poly7[58])
         );
  CFD2QXL \Poly6_reg[13]  ( .D(n9680), .CP(clk), .CD(n18342), .Q(Poly6[13]) );
  CFD2QXL \Poly15_reg[30]  ( .D(n9607), .CP(clk), .CD(n18344), .Q(Poly15[30])
         );
  CFD2QXL \Poly15_reg[29]  ( .D(n9608), .CP(clk), .CD(n18345), .Q(Poly15[29])
         );
  CFD2QXL \Poly0_reg[111]  ( .D(n9466), .CP(clk), .CD(n18350), .Q(Poly0[111])
         );
  CFD2QXL \Poly0_reg[118]  ( .D(n9459), .CP(clk), .CD(n18351), .Q(Poly0[118])
         );
  CFD2QXL \Poly0_reg[115]  ( .D(n9462), .CP(clk), .CD(n18352), .Q(Poly0[115])
         );
  CFD2QXL \Poly0_reg[120]  ( .D(n9457), .CP(clk), .CD(n18352), .Q(Poly0[120])
         );
  CFD2QXL \Poly0_reg[106]  ( .D(n9471), .CP(clk), .CD(n18353), .Q(Poly0[106])
         );
  CFD2QXL \Poly0_reg[107]  ( .D(n9470), .CP(clk), .CD(n18356), .Q(Poly0[107])
         );
  CFD2QXL \Poly1_reg[22]  ( .D(n9335), .CP(clk), .CD(n18358), .Q(Poly1[22]) );
  CFD2QXL \Poly1_reg[27]  ( .D(n9330), .CP(clk), .CD(n18360), .Q(Poly1[27]) );
  CFD2QXL \Poly1_reg[26]  ( .D(n9331), .CP(clk), .CD(n18361), .Q(Poly1[26]) );
  CFD2QXL \Poly1_reg[24]  ( .D(n9333), .CP(clk), .CD(n18363), .Q(Poly1[24]) );
  CFD2QXL \Poly1_reg[21]  ( .D(n9336), .CP(clk), .CD(n18366), .Q(Poly1[21]) );
  CFD2QXL \Poly1_reg[30]  ( .D(n9327), .CP(clk), .CD(n18370), .Q(Poly1[30]) );
  CFD2QXL \Poly1_reg[29]  ( .D(n9328), .CP(clk), .CD(n18371), .Q(Poly1[29]) );
  CFD2QXL \Poly1_reg[28]  ( .D(n9329), .CP(clk), .CD(n18374), .Q(Poly1[28]) );
  CFD2QXL \Poly1_reg[160]  ( .D(n9197), .CP(clk), .CD(n18375), .Q(Poly1[160])
         );
  CFD2QXL \Poly3_reg[36]  ( .D(n8904), .CP(clk), .CD(n18384), .Q(Poly3[36]) );
  CFD2QXL \Poly1_reg[6]  ( .D(n9351), .CP(clk), .CD(n18374), .Q(
        poly1_shifted[17]) );
  CFD2QXL \Poly15_reg[22]  ( .D(n9615), .CP(clk), .CD(n18346), .Q(Poly15[22])
         );
  CFD2QXL \Poly15_reg[25]  ( .D(n9612), .CP(clk), .CD(n18256), .Q(Poly15[25])
         );
  CFD2QXL \Poly5_reg[89]  ( .D(n11437), .CP(clk), .CD(n18257), .Q(Poly5[89])
         );
  CFD2QXL \Poly4_reg[28]  ( .D(n8828), .CP(clk), .CD(n18256), .Q(Poly4[28]) );
  CFD2QXL \Poly4_reg[0]  ( .D(n8856), .CP(clk), .CD(n18384), .Q(
        poly4_shifted[17]) );
  CFD2QXL \Poly0_reg[72]  ( .D(n9505), .CP(clk), .CD(n18347), .Q(
        poly0_shifted[90]) );
  CFD2QXL \Poly0_reg[198]  ( .D(n9379), .CP(clk), .CD(n18347), .Q(
        poly0_shifted[216]) );
  CFD2QXL \Poly0_reg[192]  ( .D(n9385), .CP(clk), .CD(n18348), .Q(
        poly0_shifted[210]) );
  CFD2QXL \Poly0_reg[196]  ( .D(n9381), .CP(clk), .CD(n18349), .Q(
        poly0_shifted[214]) );
  CFD2QXL \Poly0_reg[75]  ( .D(n9502), .CP(clk), .CD(n18349), .Q(
        poly0_shifted[93]) );
  CFD2QXL \Poly0_reg[77]  ( .D(n9500), .CP(clk), .CD(n18350), .Q(
        poly0_shifted[95]) );
  CFD2QXL \Poly0_reg[64]  ( .D(n9513), .CP(clk), .CD(n18351), .Q(
        poly0_shifted[82]) );
  CFD2QXL \Poly0_reg[66]  ( .D(n9511), .CP(clk), .CD(n18352), .Q(
        poly0_shifted[84]) );
  CFD2QXL \Poly0_reg[193]  ( .D(n9384), .CP(clk), .CD(n18352), .Q(
        poly0_shifted[211]) );
  CFD2QXL \Poly0_reg[68]  ( .D(n9509), .CP(clk), .CD(n18353), .Q(
        poly0_shifted[86]) );
  CFD2QXL \Poly0_reg[195]  ( .D(n9382), .CP(clk), .CD(n18353), .Q(
        poly0_shifted[213]) );
  CFD2QXL \Poly0_reg[65]  ( .D(n9512), .CP(clk), .CD(n18353), .Q(
        poly0_shifted[83]) );
  CFD2QXL \Poly0_reg[70]  ( .D(n9507), .CP(clk), .CD(n18353), .Q(
        poly0_shifted[88]) );
  CFD2QXL \Poly0_reg[67]  ( .D(n9510), .CP(clk), .CD(n18354), .Q(
        poly0_shifted[85]) );
  CFD2QXL \Poly0_reg[74]  ( .D(n9503), .CP(clk), .CD(n18355), .Q(
        poly0_shifted[92]) );
  CFD2QXL \Poly0_reg[201]  ( .D(n9376), .CP(clk), .CD(n18356), .Q(
        poly0_shifted[219]) );
  CFD2QXL \Poly0_reg[76]  ( .D(n9501), .CP(clk), .CD(n18356), .Q(
        poly0_shifted[94]) );
  CFD2QXL \Poly0_reg[73]  ( .D(n9504), .CP(clk), .CD(n18357), .Q(
        poly0_shifted[91]) );
  CFD2QXL \Poly1_reg[0]  ( .D(n9357), .CP(clk), .CD(n18358), .Q(
        poly1_shifted[11]) );
  CFD2QXL \Poly1_reg[11]  ( .D(n9346), .CP(clk), .CD(n18358), .Q(
        poly1_shifted[22]) );
  CFD2QXL \Poly1_reg[5]  ( .D(n9352), .CP(clk), .CD(n18360), .Q(
        poly1_shifted[16]) );
  CFD2QXL \Poly1_reg[16]  ( .D(n9341), .CP(clk), .CD(n18360), .Q(
        poly1_shifted[27]) );
  CFD2QXL \Poly1_reg[4]  ( .D(n9353), .CP(clk), .CD(n18360), .Q(
        poly1_shifted[15]) );
  CFD2QXL \Poly1_reg[15]  ( .D(n9342), .CP(clk), .CD(n18361), .Q(
        poly1_shifted[26]) );
  CFD2QXL \Poly1_reg[3]  ( .D(n9354), .CP(clk), .CD(n18361), .Q(
        poly1_shifted[14]) );
  CFD2QXL \Poly1_reg[14]  ( .D(n9343), .CP(clk), .CD(n18361), .Q(
        poly1_shifted[25]) );
  CFD2QXL \Poly1_reg[2]  ( .D(n9355), .CP(clk), .CD(n18363), .Q(
        poly1_shifted[13]) );
  CFD2QXL \Poly1_reg[13]  ( .D(n9344), .CP(clk), .CD(n18363), .Q(
        poly1_shifted[24]) );
  CFD2QXL \Poly1_reg[1]  ( .D(n9356), .CP(clk), .CD(n18364), .Q(
        poly1_shifted[12]) );
  CFD2QXL \Poly1_reg[12]  ( .D(n9345), .CP(clk), .CD(n18365), .Q(
        poly1_shifted[23]) );
  CFD2QXL \Poly1_reg[10]  ( .D(n9347), .CP(clk), .CD(n18366), .Q(
        poly1_shifted[21]) );
  CFD2QXL \Poly1_reg[9]  ( .D(n9348), .CP(clk), .CD(n18368), .Q(
        poly1_shifted[20]) );
  CFD2QXL \Poly1_reg[8]  ( .D(n9349), .CP(clk), .CD(n18370), .Q(
        poly1_shifted[19]) );
  CFD2QXL \Poly1_reg[19]  ( .D(n9338), .CP(clk), .CD(n18370), .Q(
        poly1_shifted[30]) );
  CFD2QXL \Poly1_reg[7]  ( .D(n9350), .CP(clk), .CD(n18371), .Q(
        poly1_shifted[18]) );
  CFD2QXL \Poly1_reg[18]  ( .D(n9339), .CP(clk), .CD(n18371), .Q(
        poly1_shifted[29]) );
  CFD2QXL \Poly1_reg[17]  ( .D(n9340), .CP(clk), .CD(n18374), .Q(
        poly1_shifted[28]) );
  CFD2QXL \Poly5_reg[105]  ( .D(n11421), .CP(clk), .CD(n18259), .Q(
        poly5_shifted[119]) );
  CFD2QXL \Poly5_reg[64]  ( .D(n11462), .CP(clk), .CD(n18259), .Q(
        poly5_shifted[78]) );
  CFD2QXL \Poly5_reg[109]  ( .D(n11417), .CP(clk), .CD(n18257), .Q(
        poly5_shifted[123]) );
  CFD2QXL \Poly5_reg[32]  ( .D(n11494), .CP(clk), .CD(n18257), .Q(
        poly5_shifted[46]) );
  CFD2QXL \Poly5_reg[60]  ( .D(n11466), .CP(clk), .CD(n18257), .Q(
        poly5_shifted[74]) );
  CFD2QXL \Poly8_reg[42]  ( .D(n11359), .CP(clk), .CD(n18257), .Q(
        poly8_shifted[56]) );
  CFD2QXL \Poly8_reg[56]  ( .D(n11345), .CP(clk), .CD(n18257), .Q(
        poly8_shifted[70]) );
  CFD2QXL \Poly8_reg[29]  ( .D(n11372), .CP(clk), .CD(n18257), .Q(
        poly8_shifted[43]) );
  CFD2QXL \Poly8_reg[27]  ( .D(n11374), .CP(clk), .CD(n18261), .Q(
        poly8_shifted[41]) );
  CFD2QXL \Poly8_reg[55]  ( .D(n11346), .CP(clk), .CD(n18261), .Q(
        poly8_shifted[69]) );
  CFD2QXL \Poly8_reg[40]  ( .D(n11361), .CP(clk), .CD(n18261), .Q(
        poly8_shifted[54]) );
  CFD2QXL \Poly8_reg[53]  ( .D(n11348), .CP(clk), .CD(n18261), .Q(
        poly8_shifted[67]) );
  CFD2QXL \Poly8_reg[66]  ( .D(n11335), .CP(clk), .CD(n18257), .Q(
        poly8_shifted[80]) );
  CFD2QXL \Poly8_reg[65]  ( .D(n11336), .CP(clk), .CD(n18257), .Q(
        poly8_shifted[79]) );
  CFD2QXL \Poly8_reg[19]  ( .D(n11382), .CP(clk), .CD(n18257), .Q(
        poly8_shifted[33]) );
  CFD2QXL \Poly8_reg[35]  ( .D(n11366), .CP(clk), .CD(n18257), .Q(
        poly8_shifted[49]) );
  CFD2QXL \Poly8_reg[49]  ( .D(n11352), .CP(clk), .CD(n18257), .Q(
        poly8_shifted[63]) );
  CFD2QXL \Poly8_reg[46]  ( .D(n11355), .CP(clk), .CD(n18257), .Q(
        poly8_shifted[60]) );
  CFD2QXL \Poly8_reg[60]  ( .D(n11341), .CP(clk), .CD(n18257), .Q(
        poly8_shifted[74]) );
  CFD2QXL \Poly8_reg[48]  ( .D(n11353), .CP(clk), .CD(n18257), .Q(
        poly8_shifted[62]) );
  CFD2QXL \Poly8_reg[62]  ( .D(n11339), .CP(clk), .CD(n18257), .Q(
        poly8_shifted[76]) );
  CFD2QXL \Poly9_reg[0]  ( .D(n11305), .CP(clk), .CD(n18257), .Q(
        poly9_shifted[11]) );
  CFD2QXL \Poly9_reg[55]  ( .D(n11250), .CP(clk), .CD(n18257), .Q(
        poly9_shifted[66]) );
  CFD2QXL \Poly9_reg[66]  ( .D(n11239), .CP(clk), .CD(n18257), .Q(
        poly9_shifted[77]) );
  CFD2QXL \Poly9_reg[77]  ( .D(n11228), .CP(clk), .CD(n18257), .Q(
        poly9_shifted[88]) );
  CFD2QXL \Poly9_reg[5]  ( .D(n11300), .CP(clk), .CD(n18257), .Q(
        poly9_shifted[16]) );
  CFD2QXL \Poly9_reg[6]  ( .D(n11299), .CP(clk), .CD(n18257), .Q(
        poly9_shifted[17]) );
  CFD2QXL \Poly9_reg[102]  ( .D(n11203), .CP(clk), .CD(n18257), .Q(
        poly9_shifted[113]) );
  CFD2QXL \Poly9_reg[103]  ( .D(n11202), .CP(clk), .CD(n18257), .Q(
        poly9_shifted[114]) );
  CFD2QXL \Poly9_reg[9]  ( .D(n11296), .CP(clk), .CD(n18257), .Q(
        poly9_shifted[20]) );
  CFD2QXL \Poly9_reg[104]  ( .D(n11201), .CP(clk), .CD(n18257), .Q(
        poly9_shifted[115]) );
  CFD2QXL \Poly9_reg[10]  ( .D(n11295), .CP(clk), .CD(n18257), .Q(
        poly9_shifted[21]) );
  CFD2QXL \Poly9_reg[43]  ( .D(n11262), .CP(clk), .CD(n18257), .Q(
        poly9_shifted[54]) );
  CFD2QXL \Poly9_reg[54]  ( .D(n11251), .CP(clk), .CD(n18257), .Q(
        poly9_shifted[65]) );
  CFD2QXL \Poly9_reg[1]  ( .D(n11304), .CP(clk), .CD(n18257), .Q(
        poly9_shifted[12]) );
  CFD2QXL \Poly9_reg[12]  ( .D(n11293), .CP(clk), .CD(n18257), .Q(
        poly9_shifted[23]) );
  CFD2QXL \Poly9_reg[45]  ( .D(n11260), .CP(clk), .CD(n18257), .Q(
        poly9_shifted[56]) );
  CFD2QXL \Poly9_reg[2]  ( .D(n11303), .CP(clk), .CD(n18257), .Q(
        poly9_shifted[13]) );
  CFD2QXL \Poly9_reg[46]  ( .D(n11259), .CP(clk), .CD(n18257), .Q(
        poly9_shifted[57]) );
  CFD2QXL \Poly9_reg[29]  ( .D(n11276), .CP(clk), .CD(n18257), .Q(
        poly9_shifted[40]) );
  CFD2QXL \Poly9_reg[51]  ( .D(n11254), .CP(clk), .CD(n18257), .Q(
        poly9_shifted[62]) );
  CFD2QXL \Poly9_reg[62]  ( .D(n11243), .CP(clk), .CD(n18257), .Q(
        poly9_shifted[73]) );
  CFD2QXL \Poly9_reg[73]  ( .D(n11232), .CP(clk), .CD(n18257), .Q(
        poly9_shifted[84]) );
  CFD2QXL \Poly9_reg[36]  ( .D(n11269), .CP(clk), .CD(n18257), .Q(
        poly9_shifted[47]) );
  CFD2QXL \Poly9_reg[58]  ( .D(n11247), .CP(clk), .CD(n18257), .Q(
        poly9_shifted[69]) );
  CFD2QXL \Poly9_reg[27]  ( .D(n11278), .CP(clk), .CD(n18257), .Q(
        poly9_shifted[38]) );
  CFD2QXL \Poly9_reg[71]  ( .D(n11234), .CP(clk), .CD(n18257), .Q(
        poly9_shifted[82]) );
  CFD2QXL \Poly9_reg[82]  ( .D(n11223), .CP(clk), .CD(n18257), .Q(
        poly9_shifted[93]) );
  CFD2QXL \Poly9_reg[30]  ( .D(n11275), .CP(clk), .CD(n18257), .Q(
        poly9_shifted[41]) );
  CFD2QXL \Poly9_reg[63]  ( .D(n11242), .CP(clk), .CD(n18257), .Q(
        poly9_shifted[74]) );
  CFD2QXL \Poly9_reg[74]  ( .D(n11231), .CP(clk), .CD(n18257), .Q(
        poly9_shifted[85]) );
  CFD2QXL \Poly9_reg[4]  ( .D(n11301), .CP(clk), .CD(n18257), .Q(
        poly9_shifted[15]) );
  CFD2QXL \Poly9_reg[59]  ( .D(n11246), .CP(clk), .CD(n18257), .Q(
        poly9_shifted[70]) );
  CFD2QXL \Poly9_reg[70]  ( .D(n11235), .CP(clk), .CD(n18257), .Q(
        poly9_shifted[81]) );
  CFD2QXL \Poly9_reg[81]  ( .D(n11224), .CP(clk), .CD(n18257), .Q(
        poly9_shifted[92]) );
  CFD2QXL \Poly9_reg[39]  ( .D(n11266), .CP(clk), .CD(n18257), .Q(
        poly9_shifted[50]) );
  CFD2QXL \Poly9_reg[50]  ( .D(n11255), .CP(clk), .CD(n18257), .Q(
        poly9_shifted[61]) );
  CFD2QXL \Poly9_reg[61]  ( .D(n11244), .CP(clk), .CD(n18257), .Q(
        poly9_shifted[72]) );
  CFD2QXL \Poly9_reg[72]  ( .D(n11233), .CP(clk), .CD(n18257), .Q(
        poly9_shifted[83]) );
  CFD2QXL \Poly9_reg[83]  ( .D(n11222), .CP(clk), .CD(n18257), .Q(
        poly9_shifted[94]) );
  CFD2QXL \Poly9_reg[64]  ( .D(n11241), .CP(clk), .CD(n18257), .Q(
        poly9_shifted[75]) );
  CFD2QXL \Poly11_reg[15]  ( .D(n11174), .CP(clk), .CD(n18257), .Q(
        poly11_shifted[30]) );
  CFD2QXL \Poly11_reg[3]  ( .D(n11186), .CP(clk), .CD(n18257), .Q(
        poly11_shifted[18]) );
  CFD2QXL \Poly11_reg[10]  ( .D(n11179), .CP(clk), .CD(n18257), .Q(
        poly11_shifted[25]) );
  CFD2QXL \Poly11_reg[2]  ( .D(n11187), .CP(clk), .CD(n18257), .Q(
        poly11_shifted[17]) );
  CFD2QXL \Poly11_reg[1]  ( .D(n11188), .CP(clk), .CD(n18257), .Q(
        poly11_shifted[16]) );
  CFD2QXL \Poly11_reg[16]  ( .D(n11173), .CP(clk), .CD(n18257), .Q(
        poly11_shifted[31]) );
  CFD2QXL \Poly11_reg[13]  ( .D(n11176), .CP(clk), .CD(n18257), .Q(
        poly11_shifted[28]) );
  CFD2QXL \Poly11_reg[5]  ( .D(n11184), .CP(clk), .CD(n18257), .Q(
        poly11_shifted[20]) );
  CFD2QXL \Poly13_reg[0]  ( .D(n11060), .CP(clk), .CD(n18264), .Q(
        poly13_shifted[14]) );
  CFD2QXL \Poly13_reg[42]  ( .D(n11018), .CP(clk), .CD(n18264), .Q(
        poly13_shifted[56]) );
  CFD2QXL \Poly13_reg[56]  ( .D(n11004), .CP(clk), .CD(n18264), .Q(
        poly13_shifted[70]) );
  CFD2QXL \Poly13_reg[70]  ( .D(n10990), .CP(clk), .CD(n18264), .Q(
        poly13_shifted[84]) );
  CFD2QXL \Poly13_reg[84]  ( .D(n10976), .CP(clk), .CD(n18264), .Q(
        poly13_shifted[98]) );
  CFD2QXL \Poly13_reg[98]  ( .D(n10962), .CP(clk), .CD(n18264), .Q(
        poly13_shifted[112]) );
  CFD2QXL \Poly13_reg[112]  ( .D(n10948), .CP(clk), .CD(n18264), .Q(
        poly13_shifted[126]) );
  CFD2QXL \Poly13_reg[126]  ( .D(n10934), .CP(clk), .CD(n18264), .Q(
        poly13_shifted[140]) );
  CFD2QXL \Poly13_reg[196]  ( .D(n10864), .CP(clk), .CD(n18265), .Q(
        poly13_shifted[210]) );
  CFD2QXL \Poly13_reg[210]  ( .D(n10850), .CP(clk), .CD(n18265), .Q(
        poly13_shifted[224]) );
  CFD2QXL \Poly13_reg[224]  ( .D(n10836), .CP(clk), .CD(n18265), .Q(
        poly13_shifted[238]) );
  CFD2QXL \Poly13_reg[238]  ( .D(n10822), .CP(clk), .CD(n18265), .Q(
        poly13_shifted[252]) );
  CFD2QXL \Poly13_reg[252]  ( .D(n10808), .CP(clk), .CD(n18265), .Q(
        poly13_shifted[266]) );
  CFD2QXL \Poly13_reg[294]  ( .D(n10766), .CP(clk), .CD(n18265), .Q(
        poly13_shifted[308]) );
  CFD2QXL \Poly13_reg[308]  ( .D(n10752), .CP(clk), .CD(n18265), .Q(
        poly13_shifted[322]) );
  CFD2QXL \Poly13_reg[322]  ( .D(n10738), .CP(clk), .CD(n18265), .Q(
        poly13_shifted[336]) );
  CFD2QXL \Poly13_reg[336]  ( .D(n10724), .CP(clk), .CD(n18265), .Q(
        poly13_shifted[350]) );
  CFD2QXL \Poly13_reg[350]  ( .D(n10710), .CP(clk), .CD(n18265), .Q(
        poly13_shifted[364]) );
  CFD2QXL \Poly13_reg[364]  ( .D(n10696), .CP(clk), .CD(n18265), .Q(
        poly13_shifted[378]) );
  CFD2QXL \Poly13_reg[378]  ( .D(n10682), .CP(clk), .CD(n18265), .Q(
        poly13_shifted[392]) );
  CFD2QXL \Poly13_reg[420]  ( .D(n10640), .CP(clk), .CD(n18266), .Q(
        poly13_shifted[434]) );
  CFD2QXL \Poly13_reg[434]  ( .D(n10626), .CP(clk), .CD(n18266), .Q(
        poly13_shifted[448]) );
  CFD2QXL \Poly13_reg[448]  ( .D(n10612), .CP(clk), .CD(n18266), .Q(
        poly13_shifted[462]) );
  CFD2QXL \Poly13_reg[462]  ( .D(n10598), .CP(clk), .CD(n18266), .Q(
        poly13_shifted[476]) );
  CFD2QXL \Poly13_reg[476]  ( .D(n10584), .CP(clk), .CD(n18266), .Q(
        poly13_shifted[490]) );
  CFD2QXL \Poly13_reg[490]  ( .D(n10570), .CP(clk), .CD(n18266), .Q(
        poly13_shifted[504]) );
  CFD2QXL \Poly13_reg[504]  ( .D(n10556), .CP(clk), .CD(n18266), .Q(
        poly13_shifted[518]) );
  CFD2QXL \Poly13_reg[4]  ( .D(n11056), .CP(clk), .CD(n18266), .Q(
        poly13_shifted[18]) );
  CFD2QXL \Poly13_reg[46]  ( .D(n11014), .CP(clk), .CD(n18266), .Q(
        poly13_shifted[60]) );
  CFD2QXL \Poly13_reg[74]  ( .D(n10986), .CP(clk), .CD(n18266), .Q(
        poly13_shifted[88]) );
  CFD2QXL \Poly13_reg[88]  ( .D(n10972), .CP(clk), .CD(n18267), .Q(
        poly13_shifted[102]) );
  CFD2QXL \Poly13_reg[102]  ( .D(n10958), .CP(clk), .CD(n18267), .Q(
        poly13_shifted[116]) );
  CFD2QXL \Poly13_reg[116]  ( .D(n10944), .CP(clk), .CD(n18267), .Q(
        poly13_shifted[130]) );
  CFD2QXL \Poly13_reg[130]  ( .D(n10930), .CP(clk), .CD(n18267), .Q(
        poly13_shifted[144]) );
  CFD2QXL \Poly13_reg[144]  ( .D(n10916), .CP(clk), .CD(n18267), .Q(
        poly13_shifted[158]) );
  CFD2QXL \Poly13_reg[405]  ( .D(n10655), .CP(clk), .CD(n18267), .Q(
        poly13_shifted[419]) );
  CFD2QXL \Poly13_reg[419]  ( .D(n10641), .CP(clk), .CD(n18267), .Q(
        poly13_shifted[433]) );
  CFD2QXL \Poly13_reg[433]  ( .D(n10627), .CP(clk), .CD(n18267), .Q(
        poly13_shifted[447]) );
  CFD2QXL \Poly13_reg[447]  ( .D(n10613), .CP(clk), .CD(n18267), .Q(
        poly13_shifted[461]) );
  CFD2QXL \Poly13_reg[461]  ( .D(n10599), .CP(clk), .CD(n18267), .Q(
        poly13_shifted[475]) );
  CFD2QXL \Poly13_reg[475]  ( .D(n10585), .CP(clk), .CD(n18267), .Q(
        poly13_shifted[489]) );
  CFD2QXL \Poly13_reg[489]  ( .D(n10571), .CP(clk), .CD(n18267), .Q(
        poly13_shifted[503]) );
  CFD2QXL \Poly13_reg[503]  ( .D(n10557), .CP(clk), .CD(n18267), .Q(
        poly13_shifted[517]) );
  CFD2QXL \Poly13_reg[3]  ( .D(n11057), .CP(clk), .CD(n18267), .Q(
        poly13_shifted[17]) );
  CFD2QXL \Poly13_reg[17]  ( .D(n11043), .CP(clk), .CD(n18268), .Q(
        poly13_shifted[31]) );
  CFD2QXL \Poly13_reg[31]  ( .D(n11029), .CP(clk), .CD(n18268), .Q(
        poly13_shifted[45]) );
  CFD2QXL \Poly13_reg[45]  ( .D(n11015), .CP(clk), .CD(n18268), .Q(
        poly13_shifted[59]) );
  CFD2QXL \Poly13_reg[59]  ( .D(n11001), .CP(clk), .CD(n18268), .Q(
        poly13_shifted[73]) );
  CFD2QXL \Poly13_reg[73]  ( .D(n10987), .CP(clk), .CD(n18268), .Q(
        poly13_shifted[87]) );
  CFD2QXL \Poly13_reg[87]  ( .D(n10973), .CP(clk), .CD(n18268), .Q(
        poly13_shifted[101]) );
  CFD2QXL \Poly13_reg[101]  ( .D(n10959), .CP(clk), .CD(n18268), .Q(
        poly13_shifted[115]) );
  CFD2QXL \Poly13_reg[115]  ( .D(n10945), .CP(clk), .CD(n18268), .Q(
        poly13_shifted[129]) );
  CFD2QXL \Poly13_reg[129]  ( .D(n10931), .CP(clk), .CD(n18268), .Q(
        poly13_shifted[143]) );
  CFD2QXL \Poly13_reg[143]  ( .D(n10917), .CP(clk), .CD(n18268), .Q(
        poly13_shifted[157]) );
  CFD2QXL \Poly13_reg[186]  ( .D(n10874), .CP(clk), .CD(n18268), .Q(
        poly13_shifted[200]) );
  CFD2QXL \Poly13_reg[200]  ( .D(n10860), .CP(clk), .CD(n18268), .Q(
        poly13_shifted[214]) );
  CFD2QXL \Poly13_reg[214]  ( .D(n10846), .CP(clk), .CD(n18268), .Q(
        poly13_shifted[228]) );
  CFD2QXL \Poly13_reg[228]  ( .D(n10832), .CP(clk), .CD(n18268), .Q(
        poly13_shifted[242]) );
  CFD2QXL \Poly13_reg[242]  ( .D(n10818), .CP(clk), .CD(n18269), .Q(
        poly13_shifted[256]) );
  CFD2QXL \Poly13_reg[256]  ( .D(n10804), .CP(clk), .CD(n18269), .Q(
        poly13_shifted[270]) );
  CFD2QXL \Poly13_reg[404]  ( .D(n10656), .CP(clk), .CD(n18269), .Q(
        poly13_shifted[418]) );
  CFD2QXL \Poly13_reg[446]  ( .D(n10614), .CP(clk), .CD(n18269), .Q(
        poly13_shifted[460]) );
  CFD2QXL \Poly13_reg[460]  ( .D(n10600), .CP(clk), .CD(n18269), .Q(
        poly13_shifted[474]) );
  CFD2QXL \Poly13_reg[474]  ( .D(n10586), .CP(clk), .CD(n18269), .Q(
        poly13_shifted[488]) );
  CFD2QXL \Poly13_reg[488]  ( .D(n10572), .CP(clk), .CD(n18269), .Q(
        poly13_shifted[502]) );
  CFD2QXL \Poly13_reg[502]  ( .D(n10558), .CP(clk), .CD(n18269), .Q(
        poly13_shifted[516]) );
  CFD2QXL \Poly13_reg[30]  ( .D(n11030), .CP(clk), .CD(n18269), .Q(
        poly13_shifted[44]) );
  CFD2QXL \Poly13_reg[44]  ( .D(n11016), .CP(clk), .CD(n18269), .Q(
        poly13_shifted[58]) );
  CFD2QXL \Poly13_reg[58]  ( .D(n11002), .CP(clk), .CD(n18269), .Q(
        poly13_shifted[72]) );
  CFD2QXL \Poly13_reg[100]  ( .D(n10960), .CP(clk), .CD(n18257), .Q(
        poly13_shifted[114]) );
  CFD2QXL \Poly13_reg[114]  ( .D(n10946), .CP(clk), .CD(n18257), .Q(
        poly13_shifted[128]) );
  CFD2QXL \Poly13_reg[128]  ( .D(n10932), .CP(clk), .CD(n18257), .Q(
        poly13_shifted[142]) );
  CFD2QXL \Poly13_reg[142]  ( .D(n10918), .CP(clk), .CD(n18257), .Q(
        poly13_shifted[156]) );
  CFD2QXL \Poly13_reg[185]  ( .D(n10875), .CP(clk), .CD(n18257), .Q(
        poly13_shifted[199]) );
  CFD2QXL \Poly13_reg[199]  ( .D(n10861), .CP(clk), .CD(n18257), .Q(
        poly13_shifted[213]) );
  CFD2QXL \Poly13_reg[213]  ( .D(n10847), .CP(clk), .CD(n18257), .Q(
        poly13_shifted[227]) );
  CFD2QXL \Poly13_reg[227]  ( .D(n10833), .CP(clk), .CD(n18257), .Q(
        poly13_shifted[241]) );
  CFD2QXL \Poly13_reg[403]  ( .D(n10657), .CP(clk), .CD(n18257), .Q(
        poly13_shifted[417]) );
  CFD2QXL \Poly13_reg[417]  ( .D(n10643), .CP(clk), .CD(n18257), .Q(
        poly13_shifted[431]) );
  CFD2QXL \Poly13_reg[431]  ( .D(n10629), .CP(clk), .CD(n18257), .Q(
        poly13_shifted[445]) );
  CFD2QXL \Poly13_reg[445]  ( .D(n10615), .CP(clk), .CD(n18270), .Q(
        poly13_shifted[459]) );
  CFD2QXL \Poly13_reg[459]  ( .D(n10601), .CP(clk), .CD(n18270), .Q(
        poly13_shifted[473]) );
  CFD2QXL \Poly13_reg[473]  ( .D(n10587), .CP(clk), .CD(n18270), .Q(
        poly13_shifted[487]) );
  CFD2QXL \Poly13_reg[501]  ( .D(n10559), .CP(clk), .CD(n18270), .Q(
        poly13_shifted[515]) );
  CFD2QXL \Poly13_reg[15]  ( .D(n11045), .CP(clk), .CD(n18270), .Q(
        poly13_shifted[29]) );
  CFD2QXL \Poly13_reg[57]  ( .D(n11003), .CP(clk), .CD(n18270), .Q(
        poly13_shifted[71]) );
  CFD2QXL \Poly13_reg[71]  ( .D(n10989), .CP(clk), .CD(n18270), .Q(
        poly13_shifted[85]) );
  CFD2QXL \Poly13_reg[85]  ( .D(n10975), .CP(clk), .CD(n18270), .Q(
        poly13_shifted[99]) );
  CFD2QXL \Poly13_reg[99]  ( .D(n10961), .CP(clk), .CD(n18270), .Q(
        poly13_shifted[113]) );
  CFD2QXL \Poly13_reg[141]  ( .D(n10919), .CP(clk), .CD(n18270), .Q(
        poly13_shifted[155]) );
  CFD2QXL \Poly13_reg[170]  ( .D(n10890), .CP(clk), .CD(n18271), .Q(
        poly13_shifted[184]) );
  CFD2QXL \Poly13_reg[184]  ( .D(n10876), .CP(clk), .CD(n18271), .Q(
        poly13_shifted[198]) );
  CFD2QXL \Poly13_reg[198]  ( .D(n10862), .CP(clk), .CD(n18271), .Q(
        poly13_shifted[212]) );
  CFD2QXL \Poly13_reg[226]  ( .D(n10834), .CP(clk), .CD(n18271), .Q(
        poly13_shifted[240]) );
  CFD2QXL \Poly13_reg[240]  ( .D(n10820), .CP(clk), .CD(n18271), .Q(
        poly13_shifted[254]) );
  CFD2QXL \Poly13_reg[254]  ( .D(n10806), .CP(clk), .CD(n18271), .Q(
        poly13_shifted[268]) );
  CFD2QXL \Poly13_reg[298]  ( .D(n10762), .CP(clk), .CD(n18271), .Q(
        poly13_shifted[312]) );
  CFD2QXL \Poly13_reg[312]  ( .D(n10748), .CP(clk), .CD(n18271), .Q(
        poly13_shifted[326]) );
  CFD2QXL \Poly13_reg[326]  ( .D(n10734), .CP(clk), .CD(n18271), .Q(
        poly13_shifted[340]) );
  CFD2QXL \Poly13_reg[340]  ( .D(n10720), .CP(clk), .CD(n18271), .Q(
        poly13_shifted[354]) );
  CFD2QXL \Poly13_reg[354]  ( .D(n10706), .CP(clk), .CD(n18271), .Q(
        poly13_shifted[368]) );
  CFD2QXL \Poly13_reg[368]  ( .D(n10692), .CP(clk), .CD(n18272), .Q(
        poly13_shifted[382]) );
  CFD2QXL \Poly13_reg[382]  ( .D(n10678), .CP(clk), .CD(n18272), .Q(
        poly13_shifted[396]) );
  CFD2QXL \Poly13_reg[416]  ( .D(n10644), .CP(clk), .CD(n18272), .Q(
        poly13_shifted[430]) );
  CFD2QXL \Poly13_reg[430]  ( .D(n10630), .CP(clk), .CD(n18272), .Q(
        poly13_shifted[444]) );
  CFD2QXL \Poly13_reg[444]  ( .D(n10616), .CP(clk), .CD(n18272), .Q(
        poly13_shifted[458]) );
  CFD2QXL \Poly13_reg[458]  ( .D(n10602), .CP(clk), .CD(n18272), .Q(
        poly13_shifted[472]) );
  CFD2QXL \Poly13_reg[472]  ( .D(n10588), .CP(clk), .CD(n18272), .Q(
        poly13_shifted[486]) );
  CFD2QXL \Poly13_reg[486]  ( .D(n10574), .CP(clk), .CD(n18272), .Q(
        poly13_shifted[500]) );
  CFD2QXL \Poly13_reg[500]  ( .D(n10560), .CP(clk), .CD(n18272), .Q(
        poly13_shifted[514]) );
  CFD2QXL \Poly13_reg[183]  ( .D(n10877), .CP(clk), .CD(n18272), .Q(
        poly13_shifted[197]) );
  CFD2QXL \Poly13_reg[197]  ( .D(n10863), .CP(clk), .CD(n18272), .Q(
        poly13_shifted[211]) );
  CFD2QXL \Poly13_reg[225]  ( .D(n10835), .CP(clk), .CD(n18273), .Q(
        poly13_shifted[239]) );
  CFD2QXL \Poly13_reg[239]  ( .D(n10821), .CP(clk), .CD(n18273), .Q(
        poly13_shifted[253]) );
  CFD2QXL \Poly13_reg[253]  ( .D(n10807), .CP(clk), .CD(n18273), .Q(
        poly13_shifted[267]) );
  CFD2QXL \Poly13_reg[267]  ( .D(n10793), .CP(clk), .CD(n18273), .Q(
        poly13_shifted[281]) );
  CFD2QXL \Poly13_reg[283]  ( .D(n10777), .CP(clk), .CD(n18273), .Q(
        poly13_shifted[297]) );
  CFD2QXL \Poly13_reg[297]  ( .D(n10763), .CP(clk), .CD(n18273), .Q(
        poly13_shifted[311]) );
  CFD2QXL \Poly13_reg[311]  ( .D(n10749), .CP(clk), .CD(n18273), .Q(
        poly13_shifted[325]) );
  CFD2QXL \Poly13_reg[325]  ( .D(n10735), .CP(clk), .CD(n18273), .Q(
        poly13_shifted[339]) );
  CFD2QXL \Poly13_reg[339]  ( .D(n10721), .CP(clk), .CD(n18273), .Q(
        poly13_shifted[353]) );
  CFD2QXL \Poly13_reg[353]  ( .D(n10707), .CP(clk), .CD(n18273), .Q(
        poly13_shifted[367]) );
  CFD2QXL \Poly13_reg[367]  ( .D(n10693), .CP(clk), .CD(n18273), .Q(
        poly13_shifted[381]) );
  CFD2QXL \Poly13_reg[381]  ( .D(n10679), .CP(clk), .CD(n18273), .Q(
        poly13_shifted[395]) );
  CFD2QXL \Poly13_reg[415]  ( .D(n10645), .CP(clk), .CD(n18273), .Q(
        poly13_shifted[429]) );
  CFD2QXL \Poly13_reg[429]  ( .D(n10631), .CP(clk), .CD(n18274), .Q(
        poly13_shifted[443]) );
  CFD2QXL \Poly13_reg[457]  ( .D(n10603), .CP(clk), .CD(n18274), .Q(
        poly13_shifted[471]) );
  CFD2QXL \Poly13_reg[471]  ( .D(n10589), .CP(clk), .CD(n18274), .Q(
        poly13_shifted[485]) );
  CFD2QXL \Poly13_reg[485]  ( .D(n10575), .CP(clk), .CD(n18274), .Q(
        poly13_shifted[499]) );
  CFD2QXL \Poly13_reg[499]  ( .D(n10561), .CP(clk), .CD(n18274), .Q(
        poly13_shifted[513]) );
  CFD2QXL \Poly13_reg[513]  ( .D(n10547), .CP(clk), .CD(n18274), .Q(
        poly13_shifted[527]) );
  CFD2QXL \Poly13_reg[55]  ( .D(n11005), .CP(clk), .CD(n18274), .Q(
        poly13_shifted[69]) );
  CFD2QXL \Poly13_reg[69]  ( .D(n10991), .CP(clk), .CD(n18274), .Q(
        poly13_shifted[83]) );
  CFD2QXL \Poly13_reg[83]  ( .D(n10977), .CP(clk), .CD(n18274), .Q(
        poly13_shifted[97]) );
  CFD2QXL \Poly13_reg[97]  ( .D(n10963), .CP(clk), .CD(n18274), .Q(
        poly13_shifted[111]) );
  CFD2QXL \Poly13_reg[111]  ( .D(n10949), .CP(clk), .CD(n18274), .Q(
        poly13_shifted[125]) );
  CFD2QXL \Poly13_reg[125]  ( .D(n10935), .CP(clk), .CD(n18275), .Q(
        poly13_shifted[139]) );
  CFD2QXL \Poly13_reg[139]  ( .D(n10921), .CP(clk), .CD(n18275), .Q(
        poly13_shifted[153]) );
  CFD2QXL \Poly13_reg[153]  ( .D(n10907), .CP(clk), .CD(n18275), .Q(
        poly13_shifted[167]) );
  CFD2QXL \Poly13_reg[310]  ( .D(n10750), .CP(clk), .CD(n18275), .Q(
        poly13_shifted[324]) );
  CFD2QXL \Poly13_reg[324]  ( .D(n10736), .CP(clk), .CD(n18275), .Q(
        poly13_shifted[338]) );
  CFD2QXL \Poly13_reg[366]  ( .D(n10694), .CP(clk), .CD(n18275), .Q(
        poly13_shifted[380]) );
  CFD2QXL \Poly13_reg[380]  ( .D(n10680), .CP(clk), .CD(n18275), .Q(
        poly13_shifted[394]) );
  CFD2QXL \Poly13_reg[414]  ( .D(n10646), .CP(clk), .CD(n18275), .Q(
        poly13_shifted[428]) );
  CFD2QXL \Poly13_reg[428]  ( .D(n10632), .CP(clk), .CD(n18275), .Q(
        poly13_shifted[442]) );
  CFD2QXL \Poly13_reg[442]  ( .D(n10618), .CP(clk), .CD(n18275), .Q(
        poly13_shifted[456]) );
  CFD2QXL \Poly13_reg[456]  ( .D(n10604), .CP(clk), .CD(n18275), .Q(
        poly13_shifted[470]) );
  CFD2QXL \Poly13_reg[470]  ( .D(n10590), .CP(clk), .CD(n18275), .Q(
        poly13_shifted[484]) );
  CFD2QXL \Poly13_reg[484]  ( .D(n10576), .CP(clk), .CD(n18276), .Q(
        poly13_shifted[498]) );
  CFD2QXL \Poly13_reg[498]  ( .D(n10562), .CP(clk), .CD(n18276), .Q(
        poly13_shifted[512]) );
  CFD2QXL \Poly13_reg[512]  ( .D(n10548), .CP(clk), .CD(n18276), .Q(
        poly13_shifted[526]) );
  CFD2QXL \Poly13_reg[12]  ( .D(n11048), .CP(clk), .CD(n18276), .Q(
        poly13_shifted[26]) );
  CFD2QXL \Poly13_reg[26]  ( .D(n11034), .CP(clk), .CD(n18276), .Q(
        poly13_shifted[40]) );
  CFD2QXL \Poly13_reg[40]  ( .D(n11020), .CP(clk), .CD(n18276), .Q(
        poly13_shifted[54]) );
  CFD2QXL \Poly13_reg[54]  ( .D(n11006), .CP(clk), .CD(n18276), .Q(
        poly13_shifted[68]) );
  CFD2QXL \Poly13_reg[68]  ( .D(n10992), .CP(clk), .CD(n18276), .Q(
        poly13_shifted[82]) );
  CFD2QXL \Poly13_reg[82]  ( .D(n10978), .CP(clk), .CD(n18276), .Q(
        poly13_shifted[96]) );
  CFD2QXL \Poly13_reg[124]  ( .D(n10936), .CP(clk), .CD(n18276), .Q(
        poly13_shifted[138]) );
  CFD2QXL \Poly13_reg[138]  ( .D(n10922), .CP(clk), .CD(n18276), .Q(
        poly13_shifted[152]) );
  CFD2QXL \Poly13_reg[152]  ( .D(n10908), .CP(clk), .CD(n18276), .Q(
        poly13_shifted[166]) );
  CFD2QXL \Poly13_reg[181]  ( .D(n10879), .CP(clk), .CD(n18276), .Q(
        poly13_shifted[195]) );
  CFD2QXL \Poly13_reg[195]  ( .D(n10865), .CP(clk), .CD(n18255), .Q(
        poly13_shifted[209]) );
  CFD2QXL \Poly13_reg[209]  ( .D(n10851), .CP(clk), .CD(n18255), .Q(
        poly13_shifted[223]) );
  CFD2QXL \Poly13_reg[223]  ( .D(n10837), .CP(clk), .CD(n18255), .Q(
        poly13_shifted[237]) );
  CFD2QXL \Poly13_reg[237]  ( .D(n10823), .CP(clk), .CD(n18255), .Q(
        poly13_shifted[251]) );
  CFD2QXL \Poly13_reg[251]  ( .D(n10809), .CP(clk), .CD(n18255), .Q(
        poly13_shifted[265]) );
  CFD2QXL \Poly13_reg[265]  ( .D(n10795), .CP(clk), .CD(n18255), .Q(
        poly13_shifted[279]) );
  CFD2QXL \Poly13_reg[309]  ( .D(n10751), .CP(clk), .CD(n18255), .Q(
        poly13_shifted[323]) );
  CFD2QXL \Poly13_reg[323]  ( .D(n10737), .CP(clk), .CD(n18255), .Q(
        poly13_shifted[337]) );
  CFD2QXL \Poly13_reg[337]  ( .D(n10723), .CP(clk), .CD(n18255), .Q(
        poly13_shifted[351]) );
  CFD2QXL \Poly13_reg[379]  ( .D(n10681), .CP(clk), .CD(n18255), .Q(
        poly13_shifted[393]) );
  CFD2QXL \Poly13_reg[413]  ( .D(n10647), .CP(clk), .CD(n18255), .Q(
        poly13_shifted[427]) );
  CFD2QXL \Poly13_reg[427]  ( .D(n10633), .CP(clk), .CD(n18255), .Q(
        poly13_shifted[441]) );
  CFD2QXL \Poly13_reg[441]  ( .D(n10619), .CP(clk), .CD(n18277), .Q(
        poly13_shifted[455]) );
  CFD2QXL \Poly13_reg[455]  ( .D(n10605), .CP(clk), .CD(n18277), .Q(
        poly13_shifted[469]) );
  CFD2QXL \Poly13_reg[469]  ( .D(n10591), .CP(clk), .CD(n18277), .Q(
        poly13_shifted[483]) );
  CFD2QXL \Poly13_reg[483]  ( .D(n10577), .CP(clk), .CD(n18277), .Q(
        poly13_shifted[497]) );
  CFD2QXL \Poly13_reg[511]  ( .D(n10549), .CP(clk), .CD(n18277), .Q(
        poly13_shifted[525]) );
  CFD2QXL \Poly13_reg[39]  ( .D(n11021), .CP(clk), .CD(n18277), .Q(
        poly13_shifted[53]) );
  CFD2QXL \Poly13_reg[53]  ( .D(n11007), .CP(clk), .CD(n18277), .Q(
        poly13_shifted[67]) );
  CFD2QXL \Poly13_reg[81]  ( .D(n10979), .CP(clk), .CD(n18277), .Q(
        poly13_shifted[95]) );
  CFD2QXL \Poly13_reg[95]  ( .D(n10965), .CP(clk), .CD(n18277), .Q(
        poly13_shifted[109]) );
  CFD2QXL \Poly13_reg[109]  ( .D(n10951), .CP(clk), .CD(n18277), .Q(
        poly13_shifted[123]) );
  CFD2QXL \Poly13_reg[123]  ( .D(n10937), .CP(clk), .CD(n18277), .Q(
        poly13_shifted[137]) );
  CFD2QXL \Poly13_reg[137]  ( .D(n10923), .CP(clk), .CD(n18278), .Q(
        poly13_shifted[151]) );
  CFD2QXL \Poly13_reg[180]  ( .D(n10880), .CP(clk), .CD(n18278), .Q(
        poly13_shifted[194]) );
  CFD2QXL \Poly13_reg[194]  ( .D(n10866), .CP(clk), .CD(n18278), .Q(
        poly13_shifted[208]) );
  CFD2QXL \Poly13_reg[208]  ( .D(n10852), .CP(clk), .CD(n18278), .Q(
        poly13_shifted[222]) );
  CFD2QXL \Poly13_reg[222]  ( .D(n10838), .CP(clk), .CD(n18278), .Q(
        poly13_shifted[236]) );
  CFD2QXL \Poly13_reg[236]  ( .D(n10824), .CP(clk), .CD(n18278), .Q(
        poly13_shifted[250]) );
  CFD2QXL \Poly13_reg[264]  ( .D(n10796), .CP(clk), .CD(n18278), .Q(
        poly13_shifted[278]) );
  CFD2QXL \Poly13_reg[426]  ( .D(n10634), .CP(clk), .CD(n18278), .Q(
        poly13_shifted[440]) );
  CFD2QXL \Poly13_reg[440]  ( .D(n10620), .CP(clk), .CD(n18278), .Q(
        poly13_shifted[454]) );
  CFD2QXL \Poly13_reg[454]  ( .D(n10606), .CP(clk), .CD(n18278), .Q(
        poly13_shifted[468]) );
  CFD2QXL \Poly13_reg[496]  ( .D(n10564), .CP(clk), .CD(n18279), .Q(
        poly13_shifted[510]) );
  CFD2QXL \Poly13_reg[510]  ( .D(n10550), .CP(clk), .CD(n18279), .Q(
        poly13_shifted[524]) );
  CFD2QXL \Poly13_reg[10]  ( .D(n11050), .CP(clk), .CD(n18279), .Q(
        poly13_shifted[24]) );
  CFD2QXL \Poly13_reg[24]  ( .D(n11036), .CP(clk), .CD(n18279), .Q(
        poly13_shifted[38]) );
  CFD2QXL \Poly13_reg[38]  ( .D(n11022), .CP(clk), .CD(n18279), .Q(
        poly13_shifted[52]) );
  CFD2QXL \Poly13_reg[52]  ( .D(n11008), .CP(clk), .CD(n18279), .Q(
        poly13_shifted[66]) );
  CFD2QXL \Poly13_reg[66]  ( .D(n10994), .CP(clk), .CD(n18279), .Q(
        poly13_shifted[80]) );
  CFD2QXL \Poly13_reg[80]  ( .D(n10980), .CP(clk), .CD(n18279), .Q(
        poly13_shifted[94]) );
  CFD2QXL \Poly13_reg[94]  ( .D(n10966), .CP(clk), .CD(n18279), .Q(
        poly13_shifted[108]) );
  CFD2QXL \Poly13_reg[108]  ( .D(n10952), .CP(clk), .CD(n18279), .Q(
        poly13_shifted[122]) );
  CFD2QXL \Poly13_reg[122]  ( .D(n10938), .CP(clk), .CD(n18279), .Q(
        poly13_shifted[136]) );
  CFD2QXL \Poly13_reg[136]  ( .D(n10924), .CP(clk), .CD(n18279), .Q(
        poly13_shifted[150]) );
  CFD2QXL \Poly13_reg[150]  ( .D(n10910), .CP(clk), .CD(n18279), .Q(
        poly13_shifted[164]) );
  CFD2QXL \Poly13_reg[179]  ( .D(n10881), .CP(clk), .CD(n18279), .Q(
        poly13_shifted[193]) );
  CFD2QXL \Poly13_reg[193]  ( .D(n10867), .CP(clk), .CD(n18280), .Q(
        poly13_shifted[207]) );
  CFD2QXL \Poly13_reg[207]  ( .D(n10853), .CP(clk), .CD(n18280), .Q(
        poly13_shifted[221]) );
  CFD2QXL \Poly13_reg[221]  ( .D(n10839), .CP(clk), .CD(n18280), .Q(
        poly13_shifted[235]) );
  CFD2QXL \Poly13_reg[235]  ( .D(n10825), .CP(clk), .CD(n18280), .Q(
        poly13_shifted[249]) );
  CFD2QXL \Poly13_reg[249]  ( .D(n10811), .CP(clk), .CD(n18280), .Q(
        poly13_shifted[263]) );
  CFD2QXL \Poly13_reg[263]  ( .D(n10797), .CP(clk), .CD(n18280), .Q(
        poly13_shifted[277]) );
  CFD2QXL \Poly13_reg[293]  ( .D(n10767), .CP(clk), .CD(n18280), .Q(
        poly13_shifted[307]) );
  CFD2QXL \Poly13_reg[307]  ( .D(n10753), .CP(clk), .CD(n18280), .Q(
        poly13_shifted[321]) );
  CFD2QXL \Poly13_reg[321]  ( .D(n10739), .CP(clk), .CD(n18280), .Q(
        poly13_shifted[335]) );
  CFD2QXL \Poly13_reg[335]  ( .D(n10725), .CP(clk), .CD(n18280), .Q(
        poly13_shifted[349]) );
  CFD2QXL \Poly13_reg[349]  ( .D(n10711), .CP(clk), .CD(n18280), .Q(
        poly13_shifted[363]) );
  CFD2QXL \Poly13_reg[363]  ( .D(n10697), .CP(clk), .CD(n18280), .Q(
        poly13_shifted[377]) );
  CFD2QXL \Poly13_reg[377]  ( .D(n10683), .CP(clk), .CD(n18280), .Q(
        poly13_shifted[391]) );
  CFD2QXL \Poly13_reg[439]  ( .D(n10621), .CP(clk), .CD(n18281), .Q(
        poly13_shifted[453]) );
  CFD2QXL \Poly13_reg[453]  ( .D(n10607), .CP(clk), .CD(n18281), .Q(
        poly13_shifted[467]) );
  CFD2QXL \Poly13_reg[467]  ( .D(n10593), .CP(clk), .CD(n18281), .Q(
        poly13_shifted[481]) );
  CFD2QXL \Poly13_reg[509]  ( .D(n10551), .CP(clk), .CD(n18281), .Q(
        poly13_shifted[523]) );
  CFD2QXL \Poly13_reg[9]  ( .D(n11051), .CP(clk), .CD(n18281), .Q(
        poly13_shifted[23]) );
  CFD2QXL \Poly13_reg[107]  ( .D(n10953), .CP(clk), .CD(n18281), .Q(
        poly13_shifted[121]) );
  CFD2QXL \Poly13_reg[121]  ( .D(n10939), .CP(clk), .CD(n18281), .Q(
        poly13_shifted[135]) );
  CFD2QXL \Poly13_reg[135]  ( .D(n10925), .CP(clk), .CD(n18281), .Q(
        poly13_shifted[149]) );
  CFD2QXL \Poly13_reg[149]  ( .D(n10911), .CP(clk), .CD(n18282), .Q(
        poly13_shifted[163]) );
  CFD2QXL \Poly13_reg[192]  ( .D(n10868), .CP(clk), .CD(n18282), .Q(
        poly13_shifted[206]) );
  CFD2QXL \Poly13_reg[220]  ( .D(n10840), .CP(clk), .CD(n18282), .Q(
        poly13_shifted[234]) );
  CFD2QXL \Poly13_reg[234]  ( .D(n10826), .CP(clk), .CD(n18282), .Q(
        poly13_shifted[248]) );
  CFD2QXL \Poly13_reg[248]  ( .D(n10812), .CP(clk), .CD(n18282), .Q(
        poly13_shifted[262]) );
  CFD2QXL \Poly13_reg[262]  ( .D(n10798), .CP(clk), .CD(n18282), .Q(
        poly13_shifted[276]) );
  CFD2QXL \Poly13_reg[292]  ( .D(n10768), .CP(clk), .CD(n18282), .Q(
        poly13_shifted[306]) );
  CFD2QXL \Poly13_reg[306]  ( .D(n10754), .CP(clk), .CD(n18282), .Q(
        poly13_shifted[320]) );
  CFD2QXL \Poly13_reg[320]  ( .D(n10740), .CP(clk), .CD(n18282), .Q(
        poly13_shifted[334]) );
  CFD2QXL \Poly13_reg[334]  ( .D(n10726), .CP(clk), .CD(n18282), .Q(
        poly13_shifted[348]) );
  CFD2QXL \Poly13_reg[348]  ( .D(n10712), .CP(clk), .CD(n18282), .Q(
        poly13_shifted[362]) );
  CFD2QXL \Poly13_reg[362]  ( .D(n10698), .CP(clk), .CD(n18282), .Q(
        poly13_shifted[376]) );
  CFD2QXL \Poly13_reg[424]  ( .D(n10636), .CP(clk), .CD(n18283), .Q(
        poly13_shifted[438]) );
  CFD2QXL \Poly13_reg[438]  ( .D(n10622), .CP(clk), .CD(n18283), .Q(
        poly13_shifted[452]) );
  CFD2QXL \Poly13_reg[452]  ( .D(n10608), .CP(clk), .CD(n18283), .Q(
        poly13_shifted[466]) );
  CFD2QXL \Poly13_reg[466]  ( .D(n10594), .CP(clk), .CD(n18283), .Q(
        poly13_shifted[480]) );
  CFD2QXL \Poly13_reg[480]  ( .D(n10580), .CP(clk), .CD(n18283), .Q(
        poly13_shifted[494]) );
  CFD2QXL \Poly13_reg[494]  ( .D(n10566), .CP(clk), .CD(n18283), .Q(
        poly13_shifted[508]) );
  CFD2QXL \Poly13_reg[508]  ( .D(n10552), .CP(clk), .CD(n18283), .Q(
        poly13_shifted[522]) );
  CFD2QXL \Poly13_reg[8]  ( .D(n11052), .CP(clk), .CD(n18283), .Q(
        poly13_shifted[22]) );
  CFD2QXL \Poly13_reg[22]  ( .D(n11038), .CP(clk), .CD(n18283), .Q(
        poly13_shifted[36]) );
  CFD2QXL \Poly13_reg[36]  ( .D(n11024), .CP(clk), .CD(n18283), .Q(
        poly13_shifted[50]) );
  CFD2QXL \Poly13_reg[50]  ( .D(n11010), .CP(clk), .CD(n18283), .Q(
        poly13_shifted[64]) );
  CFD2QXL \Poly13_reg[64]  ( .D(n10996), .CP(clk), .CD(n18283), .Q(
        poly13_shifted[78]) );
  CFD2QXL \Poly13_reg[78]  ( .D(n10982), .CP(clk), .CD(n18255), .Q(
        poly13_shifted[92]) );
  CFD2QXL \Poly13_reg[92]  ( .D(n10968), .CP(clk), .CD(n18255), .Q(
        poly13_shifted[106]) );
  CFD2QXL \Poly13_reg[106]  ( .D(n10954), .CP(clk), .CD(n18255), .Q(
        poly13_shifted[120]) );
  CFD2QXL \Poly13_reg[120]  ( .D(n10940), .CP(clk), .CD(n18255), .Q(
        poly13_shifted[134]) );
  CFD2QXL \Poly13_reg[134]  ( .D(n10926), .CP(clk), .CD(n18255), .Q(
        poly13_shifted[148]) );
  CFD2QXL \Poly13_reg[148]  ( .D(n10912), .CP(clk), .CD(n18255), .Q(
        poly13_shifted[162]) );
  CFD2QXL \Poly13_reg[191]  ( .D(n10869), .CP(clk), .CD(n18255), .Q(
        poly13_shifted[205]) );
  CFD2QXL \Poly13_reg[205]  ( .D(n10855), .CP(clk), .CD(n18255), .Q(
        poly13_shifted[219]) );
  CFD2QXL \Poly13_reg[233]  ( .D(n10827), .CP(clk), .CD(n18255), .Q(
        poly13_shifted[247]) );
  CFD2QXL \Poly13_reg[247]  ( .D(n10813), .CP(clk), .CD(n18255), .Q(
        poly13_shifted[261]) );
  CFD2QXL \Poly13_reg[261]  ( .D(n10799), .CP(clk), .CD(n18255), .Q(
        poly13_shifted[275]) );
  CFD2QXL \Poly13_reg[305]  ( .D(n10755), .CP(clk), .CD(n18284), .Q(
        poly13_shifted[319]) );
  CFD2QXL \Poly13_reg[319]  ( .D(n10741), .CP(clk), .CD(n18284), .Q(
        poly13_shifted[333]) );
  CFD2QXL \Poly13_reg[333]  ( .D(n10727), .CP(clk), .CD(n18284), .Q(
        poly13_shifted[347]) );
  CFD2QXL \Poly13_reg[347]  ( .D(n10713), .CP(clk), .CD(n18284), .Q(
        poly13_shifted[361]) );
  CFD2QXL \Poly13_reg[361]  ( .D(n10699), .CP(clk), .CD(n18284), .Q(
        poly13_shifted[375]) );
  CFD2QXL \Poly13_reg[375]  ( .D(n10685), .CP(clk), .CD(n18284), .Q(
        poly13_shifted[389]) );
  CFD2QXL \Poly13_reg[465]  ( .D(n10595), .CP(clk), .CD(n18284), .Q(
        poly13_shifted[479]) );
  CFD2QXL \Poly13_reg[507]  ( .D(n10553), .CP(clk), .CD(n18284), .Q(
        poly13_shifted[521]) );
  CFD2QXL \Poly13_reg[7]  ( .D(n11053), .CP(clk), .CD(n18284), .Q(
        poly13_shifted[21]) );
  CFD2QXL \Poly13_reg[21]  ( .D(n11039), .CP(clk), .CD(n18285), .Q(
        poly13_shifted[35]) );
  CFD2QXL \Poly13_reg[35]  ( .D(n11025), .CP(clk), .CD(n18285), .Q(
        poly13_shifted[49]) );
  CFD2QXL \Poly13_reg[77]  ( .D(n10983), .CP(clk), .CD(n18285), .Q(
        poly13_shifted[91]) );
  CFD2QXL \Poly13_reg[91]  ( .D(n10969), .CP(clk), .CD(n18285), .Q(
        poly13_shifted[105]) );
  CFD2QXL \Poly13_reg[105]  ( .D(n10955), .CP(clk), .CD(n18285), .Q(
        poly13_shifted[119]) );
  CFD2QXL \Poly13_reg[147]  ( .D(n10913), .CP(clk), .CD(n18285), .Q(
        poly13_shifted[161]) );
  CFD2QXL \Poly13_reg[190]  ( .D(n10870), .CP(clk), .CD(n18285), .Q(
        poly13_shifted[204]) );
  CFD2QXL \Poly13_reg[204]  ( .D(n10856), .CP(clk), .CD(n18285), .Q(
        poly13_shifted[218]) );
  CFD2QXL \Poly13_reg[218]  ( .D(n10842), .CP(clk), .CD(n18285), .Q(
        poly13_shifted[232]) );
  CFD2QXL \Poly13_reg[232]  ( .D(n10828), .CP(clk), .CD(n18285), .Q(
        poly13_shifted[246]) );
  CFD2QXL \Poly13_reg[304]  ( .D(n10756), .CP(clk), .CD(n18286), .Q(
        poly13_shifted[318]) );
  CFD2QXL \Poly13_reg[318]  ( .D(n10742), .CP(clk), .CD(n18286), .Q(
        poly13_shifted[332]) );
  CFD2QXL \Poly13_reg[332]  ( .D(n10728), .CP(clk), .CD(n18286), .Q(
        poly13_shifted[346]) );
  CFD2QXL \Poly13_reg[346]  ( .D(n10714), .CP(clk), .CD(n18286), .Q(
        poly13_shifted[360]) );
  CFD2QXL \Poly13_reg[360]  ( .D(n10700), .CP(clk), .CD(n18286), .Q(
        poly13_shifted[374]) );
  CFD2QXL \Poly13_reg[374]  ( .D(n10686), .CP(clk), .CD(n18286), .Q(
        poly13_shifted[388]) );
  CFD2QXL \Poly13_reg[408]  ( .D(n10652), .CP(clk), .CD(n18286), .Q(
        poly13_shifted[422]) );
  CFD2QXL \Poly13_reg[422]  ( .D(n10638), .CP(clk), .CD(n18286), .Q(
        poly13_shifted[436]) );
  CFD2QXL \Poly13_reg[464]  ( .D(n10596), .CP(clk), .CD(n18286), .Q(
        poly13_shifted[478]) );
  CFD2QXL \Poly13_reg[478]  ( .D(n10582), .CP(clk), .CD(n18286), .Q(
        poly13_shifted[492]) );
  CFD2QXL \Poly13_reg[492]  ( .D(n10568), .CP(clk), .CD(n18286), .Q(
        poly13_shifted[506]) );
  CFD2QXL \Poly13_reg[6]  ( .D(n11054), .CP(clk), .CD(n18287), .Q(
        poly13_shifted[20]) );
  CFD2QXL \Poly13_reg[20]  ( .D(n11040), .CP(clk), .CD(n18287), .Q(
        poly13_shifted[34]) );
  CFD2QXL \Poly13_reg[34]  ( .D(n11026), .CP(clk), .CD(n18287), .Q(
        poly13_shifted[48]) );
  CFD2QXL \Poly13_reg[48]  ( .D(n11012), .CP(clk), .CD(n18287), .Q(
        poly13_shifted[62]) );
  CFD2QXL \Poly13_reg[62]  ( .D(n10998), .CP(clk), .CD(n18287), .Q(
        poly13_shifted[76]) );
  CFD2QXL \Poly13_reg[76]  ( .D(n10984), .CP(clk), .CD(n18287), .Q(
        poly13_shifted[90]) );
  CFD2QXL \Poly13_reg[90]  ( .D(n10970), .CP(clk), .CD(n18287), .Q(
        poly13_shifted[104]) );
  CFD2QXL \Poly13_reg[104]  ( .D(n10956), .CP(clk), .CD(n18287), .Q(
        poly13_shifted[118]) );
  CFD2QXL \Poly13_reg[118]  ( .D(n10942), .CP(clk), .CD(n18287), .Q(
        poly13_shifted[132]) );
  CFD2QXL \Poly13_reg[132]  ( .D(n10928), .CP(clk), .CD(n18287), .Q(
        poly13_shifted[146]) );
  CFD2QXL \Poly13_reg[146]  ( .D(n10914), .CP(clk), .CD(n18287), .Q(
        poly13_shifted[160]) );
  CFD2QXL \Poly13_reg[189]  ( .D(n10871), .CP(clk), .CD(n18287), .Q(
        poly13_shifted[203]) );
  CFD2QXL \Poly13_reg[203]  ( .D(n10857), .CP(clk), .CD(n18288), .Q(
        poly13_shifted[217]) );
  CFD2QXL \Poly13_reg[217]  ( .D(n10843), .CP(clk), .CD(n18288), .Q(
        poly13_shifted[231]) );
  CFD2QXL \Poly13_reg[231]  ( .D(n10829), .CP(clk), .CD(n18288), .Q(
        poly13_shifted[245]) );
  CFD2QXL \Poly13_reg[245]  ( .D(n10815), .CP(clk), .CD(n18288), .Q(
        poly13_shifted[259]) );
  CFD2QXL \Poly13_reg[259]  ( .D(n10801), .CP(clk), .CD(n18288), .Q(
        poly13_shifted[273]) );
  CFD2QXL \Poly13_reg[301]  ( .D(n10759), .CP(clk), .CD(n18288), .Q(
        poly13_shifted[315]) );
  CFD2QXL \Poly13_reg[315]  ( .D(n10745), .CP(clk), .CD(n18288), .Q(
        poly13_shifted[329]) );
  CFD2QXL \Poly13_reg[359]  ( .D(n10701), .CP(clk), .CD(n18289), .Q(
        poly13_shifted[373]) );
  CFD2QXL \Poly13_reg[373]  ( .D(n10687), .CP(clk), .CD(n18289), .Q(
        poly13_shifted[387]) );
  CFD2QXL \Poly13_reg[421]  ( .D(n10639), .CP(clk), .CD(n18289), .Q(
        poly13_shifted[435]) );
  CFD2QXL \Poly13_reg[435]  ( .D(n10625), .CP(clk), .CD(n18289), .Q(
        poly13_shifted[449]) );
  CFD2QXL \Poly13_reg[449]  ( .D(n10611), .CP(clk), .CD(n18289), .Q(
        poly13_shifted[463]) );
  CFD2QXL \Poly13_reg[463]  ( .D(n10597), .CP(clk), .CD(n18289), .Q(
        poly13_shifted[477]) );
  CFD2QXL \Poly13_reg[477]  ( .D(n10583), .CP(clk), .CD(n18289), .Q(
        poly13_shifted[491]) );
  CFD2QXL \Poly13_reg[491]  ( .D(n10569), .CP(clk), .CD(n18289), .Q(
        poly13_shifted[505]) );
  CFD2QXL \Poly13_reg[47]  ( .D(n11013), .CP(clk), .CD(n18257), .Q(
        poly13_shifted[61]) );
  CFD2QXL \Poly13_reg[61]  ( .D(n10999), .CP(clk), .CD(n18257), .Q(
        poly13_shifted[75]) );
  CFD2QXL \Poly13_reg[75]  ( .D(n10985), .CP(clk), .CD(n18257), .Q(
        poly13_shifted[89]) );
  CFD2QXL \Poly13_reg[89]  ( .D(n10971), .CP(clk), .CD(n18257), .Q(
        poly13_shifted[103]) );
  CFD2QXL \Poly13_reg[103]  ( .D(n10957), .CP(clk), .CD(n18257), .Q(
        poly13_shifted[117]) );
  CFD2QXL \Poly13_reg[117]  ( .D(n10943), .CP(clk), .CD(n18257), .Q(
        poly13_shifted[131]) );
  CFD2QXL \Poly13_reg[131]  ( .D(n10929), .CP(clk), .CD(n18257), .Q(
        poly13_shifted[145]) );
  CFD2QXL \Poly13_reg[145]  ( .D(n10915), .CP(clk), .CD(n18257), .Q(
        poly13_shifted[159]) );
  CFD2QXL \Poly13_reg[173]  ( .D(n10887), .CP(clk), .CD(n18257), .Q(
        poly13_shifted[187]) );
  CFD2QXL \Poly13_reg[187]  ( .D(n10873), .CP(clk), .CD(n18257), .Q(
        poly13_shifted[201]) );
  CFD2QXL \Poly13_reg[201]  ( .D(n10859), .CP(clk), .CD(n18257), .Q(
        poly13_shifted[215]) );
  CFD2QXL \Poly13_reg[215]  ( .D(n10845), .CP(clk), .CD(n18257), .Q(
        poly13_shifted[229]) );
  CFD2QXL \Poly13_reg[229]  ( .D(n10831), .CP(clk), .CD(n18290), .Q(
        poly13_shifted[243]) );
  CFD2QXL \Poly13_reg[243]  ( .D(n10817), .CP(clk), .CD(n18290), .Q(
        poly13_shifted[257]) );
  CFD2QXL \Poly13_reg[257]  ( .D(n10803), .CP(clk), .CD(n18290), .Q(
        poly13_shifted[271]) );
  CFD2QXL \Poly13_reg[285]  ( .D(n10775), .CP(clk), .CD(n18290), .Q(
        poly13_shifted[299]) );
  CFD2QXL \Poly13_reg[327]  ( .D(n10733), .CP(clk), .CD(n18290), .Q(
        poly13_shifted[341]) );
  CFD2QXL \Poly13_reg[341]  ( .D(n10719), .CP(clk), .CD(n18290), .Q(
        poly13_shifted[355]) );
  CFD2QXL \Poly13_reg[355]  ( .D(n10705), .CP(clk), .CD(n18290), .Q(
        poly13_shifted[369]) );
  CFD2QXL \Poly13_reg[369]  ( .D(n10691), .CP(clk), .CD(n18290), .Q(
        poly13_shifted[383]) );
  CFD2QXL \Poly13_reg[383]  ( .D(n10677), .CP(clk), .CD(n18290), .Q(
        poly13_shifted[397]) );
  CFD2QXL \Poly13_reg[188]  ( .D(n10872), .CP(clk), .CD(n18290), .Q(
        poly13_shifted[202]) );
  CFD2QXL \Poly13_reg[202]  ( .D(n10858), .CP(clk), .CD(n18290), .Q(
        poly13_shifted[216]) );
  CFD2QXL \Poly13_reg[216]  ( .D(n10844), .CP(clk), .CD(n18290), .Q(
        poly13_shifted[230]) );
  CFD2QXL \Poly13_reg[230]  ( .D(n10830), .CP(clk), .CD(n18291), .Q(
        poly13_shifted[244]) );
  CFD2QXL \Poly13_reg[244]  ( .D(n10816), .CP(clk), .CD(n18291), .Q(
        poly13_shifted[258]) );
  CFD2QXL \Poly13_reg[258]  ( .D(n10802), .CP(clk), .CD(n18291), .Q(
        poly13_shifted[272]) );
  CFD2QXL \Poly13_reg[286]  ( .D(n10774), .CP(clk), .CD(n18291), .Q(
        poly13_shifted[300]) );
  CFD2QXL \Poly13_reg[300]  ( .D(n10760), .CP(clk), .CD(n18291), .Q(
        poly13_shifted[314]) );
  CFD2QXL \Poly13_reg[314]  ( .D(n10746), .CP(clk), .CD(n18291), .Q(
        poly13_shifted[328]) );
  CFD2QXL \Poly13_reg[328]  ( .D(n10732), .CP(clk), .CD(n18291), .Q(
        poly13_shifted[342]) );
  CFD2QXL \Poly13_reg[342]  ( .D(n10718), .CP(clk), .CD(n18291), .Q(
        poly13_shifted[356]) );
  CFD2QXL \Poly13_reg[356]  ( .D(n10704), .CP(clk), .CD(n18291), .Q(
        poly13_shifted[370]) );
  CFD2QXL \Poly13_reg[370]  ( .D(n10690), .CP(clk), .CD(n18291), .Q(
        poly13_shifted[384]) );
  CFD2QXL \Poly13_reg[384]  ( .D(n10676), .CP(clk), .CD(n18291), .Q(
        poly13_shifted[398]) );
  CFD2QXL \Poly13_reg[302]  ( .D(n10758), .CP(clk), .CD(n18291), .Q(
        poly13_shifted[316]) );
  CFD2QXL \Poly13_reg[316]  ( .D(n10744), .CP(clk), .CD(n18291), .Q(
        poly13_shifted[330]) );
  CFD2QXL \Poly13_reg[330]  ( .D(n10730), .CP(clk), .CD(n18292), .Q(
        poly13_shifted[344]) );
  CFD2QXL \Poly13_reg[344]  ( .D(n10716), .CP(clk), .CD(n18292), .Q(
        poly13_shifted[358]) );
  CFD2QXL \Poly13_reg[358]  ( .D(n10702), .CP(clk), .CD(n18292), .Q(
        poly13_shifted[372]) );
  CFD2QXL \Poly13_reg[372]  ( .D(n10688), .CP(clk), .CD(n18292), .Q(
        poly13_shifted[386]) );
  CFD2QXL \Poly13_reg[386]  ( .D(n10674), .CP(clk), .CD(n18292), .Q(
        poly13_shifted[400]) );
  CFD2QXL \Poly12_reg[1]  ( .D(n10531), .CP(clk), .CD(n18292), .Q(
        poly12_shifted[17]) );
  CFD2QXL \Poly12_reg[100]  ( .D(n10432), .CP(clk), .CD(n18293), .Q(
        poly12_shifted[116]) );
  CFD2QXL \Poly12_reg[6]  ( .D(n10526), .CP(clk), .CD(n18295), .Q(
        poly12_shifted[22]) );
  CFD2QXL \Poly12_reg[39]  ( .D(n10493), .CP(clk), .CD(n18295), .Q(
        poly12_shifted[55]) );
  CFD2QXL \Poly12_reg[105]  ( .D(n10427), .CP(clk), .CD(n18295), .Q(
        poly12_shifted[121]) );
  CFD2QXL \Poly12_reg[10]  ( .D(n10522), .CP(clk), .CD(n18295), .Q(
        poly12_shifted[26]) );
  CFD2QXL \Poly12_reg[75]  ( .D(n10457), .CP(clk), .CD(n18296), .Q(
        poly12_shifted[91]) );
  CFD2QXL \Poly12_reg[14]  ( .D(n10518), .CP(clk), .CD(n18297), .Q(
        poly12_shifted[30]) );
  CFD2QXL \Poly14_reg[0]  ( .D(n10405), .CP(clk), .CD(n18299), .Q(
        poly14_shifted[16]) );
  CFD2QXL \Poly14_reg[16]  ( .D(n10389), .CP(clk), .CD(n18299), .Q(
        poly14_shifted[32]) );
  CFD2QXL \Poly14_reg[32]  ( .D(n10373), .CP(clk), .CD(n18299), .Q(
        poly14_shifted[48]) );
  CFD2QXL \Poly14_reg[48]  ( .D(n10357), .CP(clk), .CD(n18299), .Q(
        poly14_shifted[64]) );
  CFD2QXL \Poly14_reg[64]  ( .D(n10341), .CP(clk), .CD(n18299), .Q(
        poly14_shifted[80]) );
  CFD2QXL \Poly14_reg[80]  ( .D(n10325), .CP(clk), .CD(n18299), .Q(
        poly14_shifted[96]) );
  CFD2QXL \Poly14_reg[96]  ( .D(n10309), .CP(clk), .CD(n18254), .Q(
        poly14_shifted[112]) );
  CFD2QXL \Poly14_reg[112]  ( .D(n10293), .CP(clk), .CD(n18254), .Q(
        poly14_shifted[128]) );
  CFD2QXL \Poly14_reg[128]  ( .D(n10277), .CP(clk), .CD(n18254), .Q(
        poly14_shifted[144]) );
  CFD2QXL \Poly14_reg[144]  ( .D(n10261), .CP(clk), .CD(n18254), .Q(
        poly14_shifted[160]) );
  CFD2QXL \Poly14_reg[160]  ( .D(n10245), .CP(clk), .CD(n18254), .Q(
        poly14_shifted[176]) );
  CFD2QXL \Poly14_reg[256]  ( .D(n10149), .CP(clk), .CD(n18254), .Q(
        poly14_shifted[272]) );
  CFD2QXL \Poly14_reg[272]  ( .D(n10133), .CP(clk), .CD(n18254), .Q(
        poly14_shifted[288]) );
  CFD2QXL \Poly14_reg[3]  ( .D(n10402), .CP(clk), .CD(n18254), .Q(
        poly14_shifted[19]) );
  CFD2QXL \Poly14_reg[19]  ( .D(n10386), .CP(clk), .CD(n18254), .Q(
        poly14_shifted[35]) );
  CFD2QXL \Poly14_reg[83]  ( .D(n10322), .CP(clk), .CD(n18300), .Q(
        poly14_shifted[99]) );
  CFD2QXL \Poly14_reg[99]  ( .D(n10306), .CP(clk), .CD(n18300), .Q(
        poly14_shifted[115]) );
  CFD2QXL \Poly14_reg[115]  ( .D(n10290), .CP(clk), .CD(n18300), .Q(
        poly14_shifted[131]) );
  CFD2QXL \Poly14_reg[131]  ( .D(n10274), .CP(clk), .CD(n18300), .Q(
        poly14_shifted[147]) );
  CFD2QXL \Poly14_reg[147]  ( .D(n10258), .CP(clk), .CD(n18300), .Q(
        poly14_shifted[163]) );
  CFD2QXL \Poly14_reg[163]  ( .D(n10242), .CP(clk), .CD(n18300), .Q(
        poly14_shifted[179]) );
  CFD2QXL \Poly14_reg[250]  ( .D(n10155), .CP(clk), .CD(n18300), .Q(
        poly14_shifted[266]) );
  CFD2QXL \Poly14_reg[266]  ( .D(n10139), .CP(clk), .CD(n18300), .Q(
        poly14_shifted[282]) );
  CFD2QXL \Poly14_reg[282]  ( .D(n10123), .CP(clk), .CD(n18300), .Q(
        poly14_shifted[298]) );
  CFD2QXL \Poly14_reg[13]  ( .D(n10392), .CP(clk), .CD(n18300), .Q(
        poly14_shifted[29]) );
  CFD2QXL \Poly14_reg[29]  ( .D(n10376), .CP(clk), .CD(n18300), .Q(
        poly14_shifted[45]) );
  CFD2QXL \Poly14_reg[45]  ( .D(n10360), .CP(clk), .CD(n18301), .Q(
        poly14_shifted[61]) );
  CFD2QXL \Poly14_reg[77]  ( .D(n10328), .CP(clk), .CD(n18301), .Q(
        poly14_shifted[93]) );
  CFD2QXL \Poly14_reg[93]  ( .D(n10312), .CP(clk), .CD(n18301), .Q(
        poly14_shifted[109]) );
  CFD2QXL \Poly14_reg[125]  ( .D(n10280), .CP(clk), .CD(n18301), .Q(
        poly14_shifted[141]) );
  CFD2QXL \Poly14_reg[141]  ( .D(n10264), .CP(clk), .CD(n18301), .Q(
        poly14_shifted[157]) );
  CFD2QXL \Poly14_reg[157]  ( .D(n10248), .CP(clk), .CD(n18301), .Q(
        poly14_shifted[173]) );
  CFD2QXL \Poly14_reg[228]  ( .D(n10177), .CP(clk), .CD(n18301), .Q(
        poly14_shifted[244]) );
  CFD2QXL \Poly14_reg[244]  ( .D(n10161), .CP(clk), .CD(n18301), .Q(
        poly14_shifted[260]) );
  CFD2QXL \Poly14_reg[260]  ( .D(n10145), .CP(clk), .CD(n18301), .Q(
        poly14_shifted[276]) );
  CFD2QXL \Poly14_reg[276]  ( .D(n10129), .CP(clk), .CD(n18301), .Q(
        poly14_shifted[292]) );
  CFD2QXL \Poly14_reg[55]  ( .D(n10350), .CP(clk), .CD(n18302), .Q(
        poly14_shifted[71]) );
  CFD2QXL \Poly14_reg[71]  ( .D(n10334), .CP(clk), .CD(n18302), .Q(
        poly14_shifted[87]) );
  CFD2QXL \Poly14_reg[87]  ( .D(n10318), .CP(clk), .CD(n18302), .Q(
        poly14_shifted[103]) );
  CFD2QXL \Poly14_reg[103]  ( .D(n10302), .CP(clk), .CD(n18302), .Q(
        poly14_shifted[119]) );
  CFD2QXL \Poly14_reg[119]  ( .D(n10286), .CP(clk), .CD(n18302), .Q(
        poly14_shifted[135]) );
  CFD2QXL \Poly14_reg[135]  ( .D(n10270), .CP(clk), .CD(n18302), .Q(
        poly14_shifted[151]) );
  CFD2QXL \Poly14_reg[151]  ( .D(n10254), .CP(clk), .CD(n18302), .Q(
        poly14_shifted[167]) );
  CFD2QXL \Poly14_reg[238]  ( .D(n10167), .CP(clk), .CD(n18302), .Q(
        poly14_shifted[254]) );
  CFD2QXL \Poly14_reg[254]  ( .D(n10151), .CP(clk), .CD(n18302), .Q(
        poly14_shifted[270]) );
  CFD2QXL \Poly14_reg[270]  ( .D(n10135), .CP(clk), .CD(n18302), .Q(
        poly14_shifted[286]) );
  CFD2QXL \Poly14_reg[17]  ( .D(n10388), .CP(clk), .CD(n18302), .Q(
        poly14_shifted[33]) );
  CFD2QXL \Poly14_reg[33]  ( .D(n10372), .CP(clk), .CD(n18303), .Q(
        poly14_shifted[49]) );
  CFD2QXL \Poly14_reg[81]  ( .D(n10324), .CP(clk), .CD(n18303), .Q(
        poly14_shifted[97]) );
  CFD2QXL \Poly14_reg[97]  ( .D(n10308), .CP(clk), .CD(n18303), .Q(
        poly14_shifted[113]) );
  CFD2QXL \Poly14_reg[113]  ( .D(n10292), .CP(clk), .CD(n18303), .Q(
        poly14_shifted[129]) );
  CFD2QXL \Poly14_reg[129]  ( .D(n10276), .CP(clk), .CD(n18303), .Q(
        poly14_shifted[145]) );
  CFD2QXL \Poly14_reg[145]  ( .D(n10260), .CP(clk), .CD(n18303), .Q(
        poly14_shifted[161]) );
  CFD2QXL \Poly14_reg[91]  ( .D(n10314), .CP(clk), .CD(n18304), .Q(
        poly14_shifted[107]) );
  CFD2QXL \Poly14_reg[107]  ( .D(n10298), .CP(clk), .CD(n18304), .Q(
        poly14_shifted[123]) );
  CFD2QXL \Poly14_reg[123]  ( .D(n10282), .CP(clk), .CD(n18304), .Q(
        poly14_shifted[139]) );
  CFD2QXL \Poly14_reg[258]  ( .D(n10147), .CP(clk), .CD(n18304), .Q(
        poly14_shifted[274]) );
  CFD2QXL \Poly14_reg[274]  ( .D(n10131), .CP(clk), .CD(n18304), .Q(
        poly14_shifted[290]) );
  CFD2QXL \Poly14_reg[21]  ( .D(n10384), .CP(clk), .CD(n18304), .Q(
        poly14_shifted[37]) );
  CFD2QXL \Poly14_reg[37]  ( .D(n10368), .CP(clk), .CD(n18304), .Q(
        poly14_shifted[53]) );
  CFD2QXL \Poly14_reg[53]  ( .D(n10352), .CP(clk), .CD(n18305), .Q(
        poly14_shifted[69]) );
  CFD2QXL \Poly14_reg[69]  ( .D(n10336), .CP(clk), .CD(n18305), .Q(
        poly14_shifted[85]) );
  CFD2QXL \Poly14_reg[85]  ( .D(n10320), .CP(clk), .CD(n18305), .Q(
        poly14_shifted[101]) );
  CFD2QXL \Poly14_reg[101]  ( .D(n10304), .CP(clk), .CD(n18305), .Q(
        poly14_shifted[117]) );
  CFD2QXL \Poly14_reg[236]  ( .D(n10169), .CP(clk), .CD(n18305), .Q(
        poly14_shifted[252]) );
  CFD2QXL \Poly14_reg[252]  ( .D(n10153), .CP(clk), .CD(n18305), .Q(
        poly14_shifted[268]) );
  CFD2QXL \Poly14_reg[268]  ( .D(n10137), .CP(clk), .CD(n18305), .Q(
        poly14_shifted[284]) );
  CFD2QXL \Poly14_reg[284]  ( .D(n10121), .CP(clk), .CD(n18305), .Q(
        poly14_shifted[300]) );
  CFD2QXL \Poly14_reg[47]  ( .D(n10358), .CP(clk), .CD(n18305), .Q(
        poly14_shifted[63]) );
  CFD2QXL \Poly14_reg[63]  ( .D(n10342), .CP(clk), .CD(n18306), .Q(
        poly14_shifted[79]) );
  CFD2QXL \Poly14_reg[79]  ( .D(n10326), .CP(clk), .CD(n18306), .Q(
        poly14_shifted[95]) );
  CFD2QXL \Poly14_reg[95]  ( .D(n10310), .CP(clk), .CD(n18306), .Q(
        poly14_shifted[111]) );
  CFD2QXL \Poly14_reg[111]  ( .D(n10294), .CP(clk), .CD(n18306), .Q(
        poly14_shifted[127]) );
  CFD2QXL \Poly14_reg[127]  ( .D(n10278), .CP(clk), .CD(n18306), .Q(
        poly14_shifted[143]) );
  CFD2QXL \Poly14_reg[143]  ( .D(n10262), .CP(clk), .CD(n18306), .Q(
        poly14_shifted[159]) );
  CFD2QXL \Poly14_reg[9]  ( .D(n10396), .CP(clk), .CD(n18306), .Q(
        poly14_shifted[25]) );
  CFD2QXL \Poly14_reg[25]  ( .D(n10380), .CP(clk), .CD(n18306), .Q(
        poly14_shifted[41]) );
  CFD2QXL \Poly14_reg[41]  ( .D(n10364), .CP(clk), .CD(n18306), .Q(
        poly14_shifted[57]) );
  CFD2QXL \Poly14_reg[89]  ( .D(n10316), .CP(clk), .CD(n18307), .Q(
        poly14_shifted[105]) );
  CFD2QXL \Poly14_reg[105]  ( .D(n10300), .CP(clk), .CD(n18307), .Q(
        poly14_shifted[121]) );
  CFD2QXL \Poly14_reg[121]  ( .D(n10284), .CP(clk), .CD(n18307), .Q(
        poly14_shifted[137]) );
  CFD2QXL \Poly14_reg[137]  ( .D(n10268), .CP(clk), .CD(n18307), .Q(
        poly14_shifted[153]) );
  CFD2QXL \Poly14_reg[233]  ( .D(n10172), .CP(clk), .CD(n18307), .Q(
        poly14_shifted[249]) );
  CFD2QXL \Poly14_reg[249]  ( .D(n10156), .CP(clk), .CD(n18307), .Q(
        poly14_shifted[265]) );
  CFD2QXL \Poly14_reg[265]  ( .D(n10140), .CP(clk), .CD(n18307), .Q(
        poly14_shifted[281]) );
  CFD2QXL \Poly14_reg[12]  ( .D(n10393), .CP(clk), .CD(n18307), .Q(
        poly14_shifted[28]) );
  CFD2QXL \Poly14_reg[28]  ( .D(n10377), .CP(clk), .CD(n18307), .Q(
        poly14_shifted[44]) );
  CFD2QXL \Poly14_reg[44]  ( .D(n10361), .CP(clk), .CD(n18308), .Q(
        poly14_shifted[60]) );
  CFD2QXL \Poly14_reg[60]  ( .D(n10345), .CP(clk), .CD(n18308), .Q(
        poly14_shifted[76]) );
  CFD2QXL \Poly14_reg[76]  ( .D(n10329), .CP(clk), .CD(n18308), .Q(
        poly14_shifted[92]) );
  CFD2QXL \Poly14_reg[92]  ( .D(n10313), .CP(clk), .CD(n18308), .Q(
        poly14_shifted[108]) );
  CFD2QXL \Poly14_reg[108]  ( .D(n10297), .CP(clk), .CD(n18308), .Q(
        poly14_shifted[124]) );
  CFD2QXL \Poly14_reg[124]  ( .D(n10281), .CP(clk), .CD(n18308), .Q(
        poly14_shifted[140]) );
  CFD2QXL \Poly14_reg[140]  ( .D(n10265), .CP(clk), .CD(n18308), .Q(
        poly14_shifted[156]) );
  CFD2QXL \Poly14_reg[156]  ( .D(n10249), .CP(clk), .CD(n18308), .Q(
        poly14_shifted[172]) );
  CFD2QXL \Poly14_reg[243]  ( .D(n10162), .CP(clk), .CD(n18308), .Q(
        poly14_shifted[259]) );
  CFD2QXL \Poly14_reg[259]  ( .D(n10146), .CP(clk), .CD(n18308), .Q(
        poly14_shifted[275]) );
  CFD2QXL \Poly14_reg[275]  ( .D(n10130), .CP(clk), .CD(n18308), .Q(
        poly14_shifted[291]) );
  CFD2QXL \Poly14_reg[6]  ( .D(n10399), .CP(clk), .CD(n18309), .Q(
        poly14_shifted[22]) );
  CFD2QXL \Poly14_reg[22]  ( .D(n10383), .CP(clk), .CD(n18309), .Q(
        poly14_shifted[38]) );
  CFD2QXL \Poly14_reg[38]  ( .D(n10367), .CP(clk), .CD(n18309), .Q(
        poly14_shifted[54]) );
  CFD2QXL \Poly14_reg[54]  ( .D(n10351), .CP(clk), .CD(n18309), .Q(
        poly14_shifted[70]) );
  CFD2QXL \Poly14_reg[70]  ( .D(n10335), .CP(clk), .CD(n18309), .Q(
        poly14_shifted[86]) );
  CFD2QXL \Poly14_reg[86]  ( .D(n10319), .CP(clk), .CD(n18309), .Q(
        poly14_shifted[102]) );
  CFD2QXL \Poly14_reg[134]  ( .D(n10271), .CP(clk), .CD(n18309), .Q(
        poly14_shifted[150]) );
  CFD2QXL \Poly14_reg[150]  ( .D(n10255), .CP(clk), .CD(n18309), .Q(
        poly14_shifted[166]) );
  CFD2QXL \Poly14_reg[187]  ( .D(n10218), .CP(clk), .CD(n18309), .Q(
        poly14_shifted[203]) );
  CFD2QXL \Poly14_reg[221]  ( .D(n10184), .CP(clk), .CD(n18310), .Q(
        poly14_shifted[237]) );
  CFD2QXL \Poly14_reg[269]  ( .D(n10136), .CP(clk), .CD(n18310), .Q(
        poly14_shifted[285]) );
  CFD2QXL \Poly14_reg[181]  ( .D(n10224), .CP(clk), .CD(n18310), .Q(
        poly14_shifted[197]) );
  CFD2QXL \Poly14_reg[247]  ( .D(n10158), .CP(clk), .CD(n18310), .Q(
        poly14_shifted[263]) );
  CFD2QXL \Poly14_reg[263]  ( .D(n10142), .CP(clk), .CD(n18310), .Q(
        poly14_shifted[279]) );
  CFD2QXL \Poly14_reg[279]  ( .D(n10126), .CP(clk), .CD(n18310), .Q(
        poly14_shifted[295]) );
  CFD2QXL \Poly14_reg[26]  ( .D(n10379), .CP(clk), .CD(n18310), .Q(
        poly14_shifted[42]) );
  CFD2QXL \Poly14_reg[42]  ( .D(n10363), .CP(clk), .CD(n18311), .Q(
        poly14_shifted[58]) );
  CFD2QXL \Poly14_reg[58]  ( .D(n10347), .CP(clk), .CD(n18311), .Q(
        poly14_shifted[74]) );
  CFD2QXL \Poly14_reg[74]  ( .D(n10331), .CP(clk), .CD(n18311), .Q(
        poly14_shifted[90]) );
  CFD2QXL \Poly14_reg[90]  ( .D(n10315), .CP(clk), .CD(n18311), .Q(
        poly14_shifted[106]) );
  CFD2QXL \Poly14_reg[122]  ( .D(n10283), .CP(clk), .CD(n18311), .Q(
        poly14_shifted[138]) );
  CFD2QXL \Poly14_reg[138]  ( .D(n10267), .CP(clk), .CD(n18311), .Q(
        poly14_shifted[154]) );
  CFD2QXL \Poly14_reg[241]  ( .D(n10164), .CP(clk), .CD(n18311), .Q(
        poly14_shifted[257]) );
  CFD2QXL \Poly14_reg[257]  ( .D(n10148), .CP(clk), .CD(n18311), .Q(
        poly14_shifted[273]) );
  CFD2QXL \Poly14_reg[4]  ( .D(n10401), .CP(clk), .CD(n18312), .Q(
        poly14_shifted[20]) );
  CFD2QXL \Poly14_reg[20]  ( .D(n10385), .CP(clk), .CD(n18312), .Q(
        poly14_shifted[36]) );
  CFD2QXL \Poly14_reg[36]  ( .D(n10369), .CP(clk), .CD(n18312), .Q(
        poly14_shifted[52]) );
  CFD2QXL \Poly14_reg[68]  ( .D(n10337), .CP(clk), .CD(n18312), .Q(
        poly14_shifted[84]) );
  CFD2QXL \Poly14_reg[84]  ( .D(n10321), .CP(clk), .CD(n18312), .Q(
        poly14_shifted[100]) );
  CFD2QXL \Poly14_reg[100]  ( .D(n10305), .CP(clk), .CD(n18312), .Q(
        poly14_shifted[116]) );
  CFD2QXL \Poly14_reg[116]  ( .D(n10289), .CP(clk), .CD(n18312), .Q(
        poly14_shifted[132]) );
  CFD2QXL \Poly14_reg[132]  ( .D(n10273), .CP(clk), .CD(n18312), .Q(
        poly14_shifted[148]) );
  CFD2QXL \Poly14_reg[148]  ( .D(n10257), .CP(clk), .CD(n18312), .Q(
        poly14_shifted[164]) );
  CFD2QXL \Poly14_reg[164]  ( .D(n10241), .CP(clk), .CD(n18312), .Q(
        poly14_shifted[180]) );
  CFD2QXL \Poly14_reg[219]  ( .D(n10186), .CP(clk), .CD(n18313), .Q(
        poly14_shifted[235]) );
  CFD2QXL \Poly14_reg[235]  ( .D(n10170), .CP(clk), .CD(n18313), .Q(
        poly14_shifted[251]) );
  CFD2QXL \Poly14_reg[251]  ( .D(n10154), .CP(clk), .CD(n18313), .Q(
        poly14_shifted[267]) );
  CFD2QXL \Poly14_reg[267]  ( .D(n10138), .CP(clk), .CD(n18313), .Q(
        poly14_shifted[283]) );
  CFD2QXL \Poly14_reg[283]  ( .D(n10122), .CP(clk), .CD(n18313), .Q(
        poly14_shifted[299]) );
  CFD2QXL \Poly14_reg[14]  ( .D(n10391), .CP(clk), .CD(n18313), .Q(
        poly14_shifted[30]) );
  CFD2QXL \Poly14_reg[30]  ( .D(n10375), .CP(clk), .CD(n18313), .Q(
        poly14_shifted[46]) );
  CFD2QXL \Poly14_reg[46]  ( .D(n10359), .CP(clk), .CD(n18313), .Q(
        poly14_shifted[62]) );
  CFD2QXL \Poly14_reg[94]  ( .D(n10311), .CP(clk), .CD(n18313), .Q(
        poly14_shifted[110]) );
  CFD2QXL \Poly14_reg[110]  ( .D(n10295), .CP(clk), .CD(n18313), .Q(
        poly14_shifted[126]) );
  CFD2QXL \Poly14_reg[126]  ( .D(n10279), .CP(clk), .CD(n18313), .Q(
        poly14_shifted[142]) );
  CFD2QXL \Poly14_reg[142]  ( .D(n10263), .CP(clk), .CD(n18313), .Q(
        poly14_shifted[158]) );
  CFD2QXL \Poly14_reg[158]  ( .D(n10247), .CP(clk), .CD(n18313), .Q(
        poly14_shifted[174]) );
  CFD2QXL \Poly14_reg[245]  ( .D(n10160), .CP(clk), .CD(n18314), .Q(
        poly14_shifted[261]) );
  CFD2QXL \Poly14_reg[261]  ( .D(n10144), .CP(clk), .CD(n18314), .Q(
        poly14_shifted[277]) );
  CFD2QXL \Poly14_reg[277]  ( .D(n10128), .CP(clk), .CD(n18314), .Q(
        poly14_shifted[293]) );
  CFD2QXL \Poly14_reg[24]  ( .D(n10381), .CP(clk), .CD(n18314), .Q(
        poly14_shifted[40]) );
  CFD2QXL \Poly14_reg[40]  ( .D(n10365), .CP(clk), .CD(n18314), .Q(
        poly14_shifted[56]) );
  CFD2QXL \Poly14_reg[56]  ( .D(n10349), .CP(clk), .CD(n18314), .Q(
        poly14_shifted[72]) );
  CFD2QXL \Poly14_reg[72]  ( .D(n10333), .CP(clk), .CD(n18314), .Q(
        poly14_shifted[88]) );
  CFD2QXL \Poly14_reg[88]  ( .D(n10317), .CP(clk), .CD(n18314), .Q(
        poly14_shifted[104]) );
  CFD2QXL \Poly14_reg[104]  ( .D(n10301), .CP(clk), .CD(n18314), .Q(
        poly14_shifted[120]) );
  CFD2QXL \Poly14_reg[120]  ( .D(n10285), .CP(clk), .CD(n18314), .Q(
        poly14_shifted[136]) );
  CFD2QXL \Poly14_reg[136]  ( .D(n10269), .CP(clk), .CD(n18314), .Q(
        poly14_shifted[152]) );
  CFD2QXL \Poly14_reg[152]  ( .D(n10253), .CP(clk), .CD(n18314), .Q(
        poly14_shifted[168]) );
  CFD2QXL \Poly14_reg[189]  ( .D(n10216), .CP(clk), .CD(n18315), .Q(
        poly14_shifted[205]) );
  CFD2QXL \Poly14_reg[239]  ( .D(n10166), .CP(clk), .CD(n18315), .Q(
        poly14_shifted[255]) );
  CFD2QXL \Poly14_reg[255]  ( .D(n10150), .CP(clk), .CD(n18315), .Q(
        poly14_shifted[271]) );
  CFD2QXL \Poly14_reg[271]  ( .D(n10134), .CP(clk), .CD(n18315), .Q(
        poly14_shifted[287]) );
  CFD2QXL \Poly14_reg[2]  ( .D(n10403), .CP(clk), .CD(n18315), .Q(
        poly14_shifted[18]) );
  CFD2QXL \Poly14_reg[18]  ( .D(n10387), .CP(clk), .CD(n18315), .Q(
        poly14_shifted[34]) );
  CFD2QXL \Poly14_reg[34]  ( .D(n10371), .CP(clk), .CD(n18315), .Q(
        poly14_shifted[50]) );
  CFD2QXL \Poly14_reg[66]  ( .D(n10339), .CP(clk), .CD(n18315), .Q(
        poly14_shifted[82]) );
  CFD2QXL \Poly14_reg[82]  ( .D(n10323), .CP(clk), .CD(n18315), .Q(
        poly14_shifted[98]) );
  CFD2QXL \Poly14_reg[98]  ( .D(n10307), .CP(clk), .CD(n18315), .Q(
        poly14_shifted[114]) );
  CFD2QXL \Poly14_reg[114]  ( .D(n10291), .CP(clk), .CD(n18316), .Q(
        poly14_shifted[130]) );
  CFD2QXL \Poly14_reg[130]  ( .D(n10275), .CP(clk), .CD(n18316), .Q(
        poly14_shifted[146]) );
  CFD2QXL \Poly14_reg[146]  ( .D(n10259), .CP(clk), .CD(n18316), .Q(
        poly14_shifted[162]) );
  CFD2QXL \Poly14_reg[190]  ( .D(n10215), .CP(clk), .CD(n18316), .Q(
        poly14_shifted[206]) );
  CFD2QXL \Poly7_reg[0]  ( .D(n10104), .CP(clk), .CD(n18316), .Q(
        poly7_shifted[12]) );
  CFD2QXL \Poly7_reg[12]  ( .D(n10092), .CP(clk), .CD(n18316), .Q(
        poly7_shifted[24]) );
  CFD2QXL \Poly7_reg[72]  ( .D(n10032), .CP(clk), .CD(n18317), .Q(
        poly7_shifted[84]) );
  CFD2QXL \Poly7_reg[84]  ( .D(n10020), .CP(clk), .CD(n18317), .Q(
        poly7_shifted[96]) );
  CFD2QXL \Poly7_reg[96]  ( .D(n10008), .CP(clk), .CD(n18317), .Q(
        poly7_shifted[108]) );
  CFD2QXL \Poly7_reg[108]  ( .D(n9996), .CP(clk), .CD(n18317), .Q(
        poly7_shifted[120]) );
  CFD2QXL \Poly7_reg[216]  ( .D(n9888), .CP(clk), .CD(n18317), .Q(
        poly7_shifted[228]) );
  CFD2QXL \Poly7_reg[228]  ( .D(n9876), .CP(clk), .CD(n18317), .Q(
        poly7_shifted[240]) );
  CFD2QXL \Poly7_reg[264]  ( .D(n9840), .CP(clk), .CD(n18318), .Q(
        poly7_shifted[276]) );
  CFD2QXL \Poly7_reg[276]  ( .D(n9828), .CP(clk), .CD(n18318), .Q(
        poly7_shifted[288]) );
  CFD2QXL \Poly7_reg[288]  ( .D(n9816), .CP(clk), .CD(n18318), .Q(
        poly7_shifted[300]) );
  CFD2QXL \Poly7_reg[300]  ( .D(n9804), .CP(clk), .CD(n18318), .Q(
        poly7_shifted[312]) );
  CFD2QXL \Poly7_reg[312]  ( .D(n9792), .CP(clk), .CD(n18318), .Q(
        poly7_shifted[324]) );
  CFD2QXL \Poly7_reg[324]  ( .D(n9780), .CP(clk), .CD(n18318), .Q(
        poly7_shifted[336]) );
  CFD2QXL \Poly7_reg[336]  ( .D(n9768), .CP(clk), .CD(n18318), .Q(
        poly7_shifted[348]) );
  CFD2QXL \Poly7_reg[348]  ( .D(n9756), .CP(clk), .CD(n18318), .Q(
        poly7_shifted[360]) );
  CFD2QXL \Poly7_reg[360]  ( .D(n9744), .CP(clk), .CD(n18318), .Q(
        poly7_shifted[372]) );
  CFD2QXL \Poly7_reg[372]  ( .D(n9732), .CP(clk), .CD(n18318), .Q(
        poly7_shifted[384]) );
  CFD2QXL \Poly7_reg[384]  ( .D(n9720), .CP(clk), .CD(n18318), .Q(
        poly7_shifted[396]) );
  CFD2QXL \Poly7_reg[396]  ( .D(n9708), .CP(clk), .CD(n18318), .Q(
        poly7_shifted[408]) );
  CFD2QXL \Poly7_reg[9]  ( .D(n10095), .CP(clk), .CD(n18318), .Q(
        poly7_shifted[21]) );
  CFD2QXL \Poly7_reg[266]  ( .D(n9838), .CP(clk), .CD(n18319), .Q(
        poly7_shifted[278]) );
  CFD2QXL \Poly7_reg[302]  ( .D(n9802), .CP(clk), .CD(n18319), .Q(
        poly7_shifted[314]) );
  CFD2QXL \Poly7_reg[314]  ( .D(n9790), .CP(clk), .CD(n18319), .Q(
        poly7_shifted[326]) );
  CFD2QXL \Poly7_reg[326]  ( .D(n9778), .CP(clk), .CD(n18319), .Q(
        poly7_shifted[338]) );
  CFD2QXL \Poly7_reg[338]  ( .D(n9766), .CP(clk), .CD(n18319), .Q(
        poly7_shifted[350]) );
  CFD2QXL \Poly7_reg[350]  ( .D(n9754), .CP(clk), .CD(n18319), .Q(
        poly7_shifted[362]) );
  CFD2QXL \Poly7_reg[362]  ( .D(n9742), .CP(clk), .CD(n18319), .Q(
        poly7_shifted[374]) );
  CFD2QXL \Poly7_reg[374]  ( .D(n9730), .CP(clk), .CD(n18319), .Q(
        poly7_shifted[386]) );
  CFD2QXL \Poly7_reg[386]  ( .D(n9718), .CP(clk), .CD(n18319), .Q(
        poly7_shifted[398]) );
  CFD2QXL \Poly7_reg[268]  ( .D(n9836), .CP(clk), .CD(n18320), .Q(
        poly7_shifted[280]) );
  CFD2QXL \Poly7_reg[280]  ( .D(n9824), .CP(clk), .CD(n18320), .Q(
        poly7_shifted[292]) );
  CFD2QXL \Poly7_reg[292]  ( .D(n9812), .CP(clk), .CD(n18320), .Q(
        poly7_shifted[304]) );
  CFD2QXL \Poly7_reg[304]  ( .D(n9800), .CP(clk), .CD(n18320), .Q(
        poly7_shifted[316]) );
  CFD2QXL \Poly7_reg[316]  ( .D(n9788), .CP(clk), .CD(n18320), .Q(
        poly7_shifted[328]) );
  CFD2QXL \Poly7_reg[328]  ( .D(n9776), .CP(clk), .CD(n18320), .Q(
        poly7_shifted[340]) );
  CFD2QXL \Poly7_reg[340]  ( .D(n9764), .CP(clk), .CD(n18320), .Q(
        poly7_shifted[352]) );
  CFD2QXL \Poly7_reg[352]  ( .D(n9752), .CP(clk), .CD(n18320), .Q(
        poly7_shifted[364]) );
  CFD2QXL \Poly7_reg[364]  ( .D(n9740), .CP(clk), .CD(n18320), .Q(
        poly7_shifted[376]) );
  CFD2QXL \Poly7_reg[376]  ( .D(n9728), .CP(clk), .CD(n18320), .Q(
        poly7_shifted[388]) );
  CFD2QXL \Poly7_reg[388]  ( .D(n9716), .CP(clk), .CD(n18320), .Q(
        poly7_shifted[400]) );
  CFD2QXL \Poly7_reg[1]  ( .D(n10103), .CP(clk), .CD(n18320), .Q(
        poly7_shifted[13]) );
  CFD2QXL \Poly7_reg[13]  ( .D(n10091), .CP(clk), .CD(n18320), .Q(
        poly7_shifted[25]) );
  CFD2QXL \Poly7_reg[258]  ( .D(n9846), .CP(clk), .CD(n18321), .Q(
        poly7_shifted[270]) );
  CFD2QXL \Poly7_reg[270]  ( .D(n9834), .CP(clk), .CD(n18321), .Q(
        poly7_shifted[282]) );
  CFD2QXL \Poly7_reg[282]  ( .D(n9822), .CP(clk), .CD(n18321), .Q(
        poly7_shifted[294]) );
  CFD2QXL \Poly7_reg[294]  ( .D(n9810), .CP(clk), .CD(n18321), .Q(
        poly7_shifted[306]) );
  CFD2QXL \Poly7_reg[306]  ( .D(n9798), .CP(clk), .CD(n18321), .Q(
        poly7_shifted[318]) );
  CFD2QXL \Poly7_reg[342]  ( .D(n9762), .CP(clk), .CD(n18321), .Q(
        poly7_shifted[354]) );
  CFD2QXL \Poly7_reg[354]  ( .D(n9750), .CP(clk), .CD(n18321), .Q(
        poly7_shifted[366]) );
  CFD2QXL \Poly7_reg[366]  ( .D(n9738), .CP(clk), .CD(n18321), .Q(
        poly7_shifted[378]) );
  CFD2QXL \Poly7_reg[3]  ( .D(n10101), .CP(clk), .CD(n18321), .Q(
        poly7_shifted[15]) );
  CFD2QXL \Poly7_reg[15]  ( .D(n10089), .CP(clk), .CD(n18321), .Q(
        poly7_shifted[27]) );
  CFD2QXL \Poly7_reg[260]  ( .D(n9844), .CP(clk), .CD(n18321), .Q(
        poly7_shifted[272]) );
  CFD2QXL \Poly7_reg[272]  ( .D(n9832), .CP(clk), .CD(n18322), .Q(
        poly7_shifted[284]) );
  CFD2QXL \Poly7_reg[284]  ( .D(n9820), .CP(clk), .CD(n18322), .Q(
        poly7_shifted[296]) );
  CFD2QXL \Poly7_reg[296]  ( .D(n9808), .CP(clk), .CD(n18322), .Q(
        poly7_shifted[308]) );
  CFD2QXL \Poly7_reg[308]  ( .D(n9796), .CP(clk), .CD(n18322), .Q(
        poly7_shifted[320]) );
  CFD2QXL \Poly7_reg[332]  ( .D(n9772), .CP(clk), .CD(n18322), .Q(
        poly7_shifted[344]) );
  CFD2QXL \Poly7_reg[344]  ( .D(n9760), .CP(clk), .CD(n18322), .Q(
        poly7_shifted[356]) );
  CFD2QXL \Poly7_reg[356]  ( .D(n9748), .CP(clk), .CD(n18322), .Q(
        poly7_shifted[368]) );
  CFD2QXL \Poly7_reg[380]  ( .D(n9724), .CP(clk), .CD(n18322), .Q(
        poly7_shifted[392]) );
  CFD2QXL \Poly7_reg[392]  ( .D(n9712), .CP(clk), .CD(n18322), .Q(
        poly7_shifted[404]) );
  CFD2QXL \Poly7_reg[17]  ( .D(n10087), .CP(clk), .CD(n18322), .Q(
        poly7_shifted[29]) );
  CFD2QXL \Poly7_reg[262]  ( .D(n9842), .CP(clk), .CD(n18323), .Q(
        poly7_shifted[274]) );
  CFD2QXL \Poly7_reg[274]  ( .D(n9830), .CP(clk), .CD(n18323), .Q(
        poly7_shifted[286]) );
  CFD2QXL \Poly7_reg[286]  ( .D(n9818), .CP(clk), .CD(n18323), .Q(
        poly7_shifted[298]) );
  CFD2QXL \Poly7_reg[298]  ( .D(n9806), .CP(clk), .CD(n18323), .Q(
        poly7_shifted[310]) );
  CFD2QXL \Poly7_reg[322]  ( .D(n9782), .CP(clk), .CD(n18323), .Q(
        poly7_shifted[334]) );
  CFD2QXL \Poly7_reg[334]  ( .D(n9770), .CP(clk), .CD(n18323), .Q(
        poly7_shifted[346]) );
  CFD2QXL \Poly7_reg[346]  ( .D(n9758), .CP(clk), .CD(n18323), .Q(
        poly7_shifted[358]) );
  CFD2QXL \Poly7_reg[358]  ( .D(n9746), .CP(clk), .CD(n18323), .Q(
        poly7_shifted[370]) );
  CFD2QXL \Poly7_reg[370]  ( .D(n9734), .CP(clk), .CD(n18323), .Q(
        poly7_shifted[382]) );
  CFD2QXL \Poly7_reg[382]  ( .D(n9722), .CP(clk), .CD(n18323), .Q(
        poly7_shifted[394]) );
  CFD2QXL \Poly7_reg[394]  ( .D(n9710), .CP(clk), .CD(n18323), .Q(
        poly7_shifted[406]) );
  CFD2QXL \Poly7_reg[7]  ( .D(n10097), .CP(clk), .CD(n18323), .Q(
        poly7_shifted[19]) );
  CFD2QXL \Poly7_reg[209]  ( .D(n9895), .CP(clk), .CD(n18323), .Q(
        poly7_shifted[221]) );
  CFD2QXL \Poly7_reg[221]  ( .D(n9883), .CP(clk), .CD(n18324), .Q(
        poly7_shifted[233]) );
  CFD2QXL \Poly7_reg[245]  ( .D(n9859), .CP(clk), .CD(n18324), .Q(
        poly7_shifted[257]) );
  CFD2QXL \Poly7_reg[257]  ( .D(n9847), .CP(clk), .CD(n18324), .Q(
        poly7_shifted[269]) );
  CFD2QXL \Poly7_reg[269]  ( .D(n9835), .CP(clk), .CD(n18324), .Q(
        poly7_shifted[281]) );
  CFD2QXL \Poly7_reg[281]  ( .D(n9823), .CP(clk), .CD(n18324), .Q(
        poly7_shifted[293]) );
  CFD2QXL \Poly7_reg[293]  ( .D(n9811), .CP(clk), .CD(n18324), .Q(
        poly7_shifted[305]) );
  CFD2QXL \Poly7_reg[305]  ( .D(n9799), .CP(clk), .CD(n18324), .Q(
        poly7_shifted[317]) );
  CFD2QXL \Poly7_reg[317]  ( .D(n9787), .CP(clk), .CD(n18324), .Q(
        poly7_shifted[329]) );
  CFD2QXL \Poly7_reg[329]  ( .D(n9775), .CP(clk), .CD(n18324), .Q(
        poly7_shifted[341]) );
  CFD2QXL \Poly7_reg[341]  ( .D(n9763), .CP(clk), .CD(n18324), .Q(
        poly7_shifted[353]) );
  CFD2QXL \Poly7_reg[353]  ( .D(n9751), .CP(clk), .CD(n18324), .Q(
        poly7_shifted[365]) );
  CFD2QXL \Poly7_reg[365]  ( .D(n9739), .CP(clk), .CD(n18324), .Q(
        poly7_shifted[377]) );
  CFD2QXL \Poly7_reg[377]  ( .D(n9727), .CP(clk), .CD(n18324), .Q(
        poly7_shifted[389]) );
  CFD2QXL \Poly7_reg[389]  ( .D(n9715), .CP(clk), .CD(n18324), .Q(
        poly7_shifted[401]) );
  CFD2QXL \Poly7_reg[2]  ( .D(n10102), .CP(clk), .CD(n18325), .Q(
        poly7_shifted[14]) );
  CFD2QXL \Poly7_reg[14]  ( .D(n10090), .CP(clk), .CD(n18325), .Q(
        poly7_shifted[26]) );
  CFD2QXL \Poly7_reg[45]  ( .D(n10059), .CP(clk), .CD(n18325), .Q(
        poly7_shifted[57]) );
  CFD2QXL \Poly7_reg[81]  ( .D(n10023), .CP(clk), .CD(n18325), .Q(
        poly7_shifted[93]) );
  CFD2QXL \Poly7_reg[93]  ( .D(n10011), .CP(clk), .CD(n18325), .Q(
        poly7_shifted[105]) );
  CFD2QXL \Poly7_reg[105]  ( .D(n9999), .CP(clk), .CD(n18325), .Q(
        poly7_shifted[117]) );
  CFD2QXL \Poly7_reg[117]  ( .D(n9987), .CP(clk), .CD(n18325), .Q(
        poly7_shifted[129]) );
  CFD2QXL \Poly7_reg[129]  ( .D(n9975), .CP(clk), .CD(n18325), .Q(
        poly7_shifted[141]) );
  CFD2QXL \Poly7_reg[141]  ( .D(n9963), .CP(clk), .CD(n18325), .Q(
        poly7_shifted[153]) );
  CFD2QXL \Poly7_reg[153]  ( .D(n9951), .CP(clk), .CD(n18326), .Q(
        poly7_shifted[165]) );
  CFD2QXL \Poly7_reg[165]  ( .D(n9939), .CP(clk), .CD(n18326), .Q(
        poly7_shifted[177]) );
  CFD2QXL \Poly7_reg[177]  ( .D(n9927), .CP(clk), .CD(n18326), .Q(
        poly7_shifted[189]) );
  CFD2QXL \Poly7_reg[74]  ( .D(n10030), .CP(clk), .CD(n18326), .Q(
        poly7_shifted[86]) );
  CFD2QXL \Poly7_reg[86]  ( .D(n10018), .CP(clk), .CD(n18326), .Q(
        poly7_shifted[98]) );
  CFD2QXL \Poly7_reg[98]  ( .D(n10006), .CP(clk), .CD(n18326), .Q(
        poly7_shifted[110]) );
  CFD2QXL \Poly7_reg[110]  ( .D(n9994), .CP(clk), .CD(n18326), .Q(
        poly7_shifted[122]) );
  CFD2QXL \Poly7_reg[122]  ( .D(n9982), .CP(clk), .CD(n18326), .Q(
        poly7_shifted[134]) );
  CFD2QXL \Poly7_reg[170]  ( .D(n9934), .CP(clk), .CD(n18326), .Q(
        poly7_shifted[182]) );
  CFD2QXL \Poly7_reg[259]  ( .D(n9845), .CP(clk), .CD(n18326), .Q(
        poly7_shifted[271]) );
  CFD2QXL \Poly7_reg[271]  ( .D(n9833), .CP(clk), .CD(n18327), .Q(
        poly7_shifted[283]) );
  CFD2QXL \Poly7_reg[283]  ( .D(n9821), .CP(clk), .CD(n18327), .Q(
        poly7_shifted[295]) );
  CFD2QXL \Poly7_reg[295]  ( .D(n9809), .CP(clk), .CD(n18327), .Q(
        poly7_shifted[307]) );
  CFD2QXL \Poly7_reg[319]  ( .D(n9785), .CP(clk), .CD(n18327), .Q(
        poly7_shifted[331]) );
  CFD2QXL \Poly7_reg[331]  ( .D(n9773), .CP(clk), .CD(n18327), .Q(
        poly7_shifted[343]) );
  CFD2QXL \Poly7_reg[343]  ( .D(n9761), .CP(clk), .CD(n18327), .Q(
        poly7_shifted[355]) );
  CFD2QXL \Poly7_reg[355]  ( .D(n9749), .CP(clk), .CD(n18327), .Q(
        poly7_shifted[367]) );
  CFD2QXL \Poly7_reg[391]  ( .D(n9713), .CP(clk), .CD(n18327), .Q(
        poly7_shifted[403]) );
  CFD2QXL \Poly7_reg[4]  ( .D(n10100), .CP(clk), .CD(n18327), .Q(
        poly7_shifted[16]) );
  CFD2QXL \Poly7_reg[16]  ( .D(n10088), .CP(clk), .CD(n18327), .Q(
        poly7_shifted[28]) );
  CFD2QXL \Poly7_reg[83]  ( .D(n10021), .CP(clk), .CD(n18328), .Q(
        poly7_shifted[95]) );
  CFD2QXL \Poly7_reg[95]  ( .D(n10009), .CP(clk), .CD(n18328), .Q(
        poly7_shifted[107]) );
  CFD2QXL \Poly7_reg[107]  ( .D(n9997), .CP(clk), .CD(n18328), .Q(
        poly7_shifted[119]) );
  CFD2QXL \Poly7_reg[119]  ( .D(n9985), .CP(clk), .CD(n18328), .Q(
        poly7_shifted[131]) );
  CFD2QXL \Poly7_reg[131]  ( .D(n9973), .CP(clk), .CD(n18328), .Q(
        poly7_shifted[143]) );
  CFD2QXL \Poly7_reg[143]  ( .D(n9961), .CP(clk), .CD(n18328), .Q(
        poly7_shifted[155]) );
  CFD2QXL \Poly7_reg[155]  ( .D(n9949), .CP(clk), .CD(n18328), .Q(
        poly7_shifted[167]) );
  CFD2QXL \Poly7_reg[167]  ( .D(n9937), .CP(clk), .CD(n18328), .Q(
        poly7_shifted[179]) );
  CFD2QXL \Poly7_reg[76]  ( .D(n10028), .CP(clk), .CD(n18329), .Q(
        poly7_shifted[88]) );
  CFD2QXL \Poly7_reg[88]  ( .D(n10016), .CP(clk), .CD(n18329), .Q(
        poly7_shifted[100]) );
  CFD2QXL \Poly7_reg[100]  ( .D(n10004), .CP(clk), .CD(n18329), .Q(
        poly7_shifted[112]) );
  CFD2QXL \Poly7_reg[112]  ( .D(n9992), .CP(clk), .CD(n18329), .Q(
        poly7_shifted[124]) );
  CFD2QXL \Poly7_reg[124]  ( .D(n9980), .CP(clk), .CD(n18329), .Q(
        poly7_shifted[136]) );
  CFD2QXL \Poly7_reg[136]  ( .D(n9968), .CP(clk), .CD(n18329), .Q(
        poly7_shifted[148]) );
  CFD2QXL \Poly7_reg[148]  ( .D(n9956), .CP(clk), .CD(n18329), .Q(
        poly7_shifted[160]) );
  CFD2QXL \Poly7_reg[160]  ( .D(n9944), .CP(clk), .CD(n18329), .Q(
        poly7_shifted[172]) );
  CFD2QXL \Poly7_reg[172]  ( .D(n9932), .CP(clk), .CD(n18329), .Q(
        poly7_shifted[184]) );
  CFD2QXL \Poly7_reg[261]  ( .D(n9843), .CP(clk), .CD(n18329), .Q(
        poly7_shifted[273]) );
  CFD2QXL \Poly7_reg[273]  ( .D(n9831), .CP(clk), .CD(n18330), .Q(
        poly7_shifted[285]) );
  CFD2QXL \Poly7_reg[285]  ( .D(n9819), .CP(clk), .CD(n18330), .Q(
        poly7_shifted[297]) );
  CFD2QXL \Poly7_reg[297]  ( .D(n9807), .CP(clk), .CD(n18330), .Q(
        poly7_shifted[309]) );
  CFD2QXL \Poly7_reg[309]  ( .D(n9795), .CP(clk), .CD(n18330), .Q(
        poly7_shifted[321]) );
  CFD2QXL \Poly7_reg[321]  ( .D(n9783), .CP(clk), .CD(n18330), .Q(
        poly7_shifted[333]) );
  CFD2QXL \Poly7_reg[333]  ( .D(n9771), .CP(clk), .CD(n18330), .Q(
        poly7_shifted[345]) );
  CFD2QXL \Poly7_reg[345]  ( .D(n9759), .CP(clk), .CD(n18330), .Q(
        poly7_shifted[357]) );
  CFD2QXL \Poly7_reg[357]  ( .D(n9747), .CP(clk), .CD(n18330), .Q(
        poly7_shifted[369]) );
  CFD2QXL \Poly7_reg[369]  ( .D(n9735), .CP(clk), .CD(n18330), .Q(
        poly7_shifted[381]) );
  CFD2QXL \Poly7_reg[381]  ( .D(n9723), .CP(clk), .CD(n18330), .Q(
        poly7_shifted[393]) );
  CFD2QXL \Poly7_reg[393]  ( .D(n9711), .CP(clk), .CD(n18330), .Q(
        poly7_shifted[405]) );
  CFD2QXL \Poly7_reg[18]  ( .D(n10086), .CP(clk), .CD(n18330), .Q(
        poly7_shifted[30]) );
  CFD2QXL \Poly7_reg[61]  ( .D(n10043), .CP(clk), .CD(n18331), .Q(
        poly7_shifted[73]) );
  CFD2QXL \Poly7_reg[97]  ( .D(n10007), .CP(clk), .CD(n18331), .Q(
        poly7_shifted[109]) );
  CFD2QXL \Poly7_reg[109]  ( .D(n9995), .CP(clk), .CD(n18331), .Q(
        poly7_shifted[121]) );
  CFD2QXL \Poly7_reg[121]  ( .D(n9983), .CP(clk), .CD(n18331), .Q(
        poly7_shifted[133]) );
  CFD2QXL \Poly7_reg[133]  ( .D(n9971), .CP(clk), .CD(n18331), .Q(
        poly7_shifted[145]) );
  CFD2QXL \Poly7_reg[145]  ( .D(n9959), .CP(clk), .CD(n18331), .Q(
        poly7_shifted[157]) );
  CFD2QXL \Poly7_reg[157]  ( .D(n9947), .CP(clk), .CD(n18331), .Q(
        poly7_shifted[169]) );
  CFD2QXL \Poly7_reg[169]  ( .D(n9935), .CP(clk), .CD(n18331), .Q(
        poly7_shifted[181]) );
  CFD2QXL \Poly7_reg[78]  ( .D(n10026), .CP(clk), .CD(n18332), .Q(
        poly7_shifted[90]) );
  CFD2QXL \Poly7_reg[114]  ( .D(n9990), .CP(clk), .CD(n18332), .Q(
        poly7_shifted[126]) );
  CFD2QXL \Poly7_reg[126]  ( .D(n9978), .CP(clk), .CD(n18332), .Q(
        poly7_shifted[138]) );
  CFD2QXL \Poly7_reg[138]  ( .D(n9966), .CP(clk), .CD(n18332), .Q(
        poly7_shifted[150]) );
  CFD2QXL \Poly7_reg[150]  ( .D(n9954), .CP(clk), .CD(n18332), .Q(
        poly7_shifted[162]) );
  CFD2QXL \Poly7_reg[162]  ( .D(n9942), .CP(clk), .CD(n18332), .Q(
        poly7_shifted[174]) );
  CFD2QXL \Poly7_reg[174]  ( .D(n9930), .CP(clk), .CD(n18332), .Q(
        poly7_shifted[186]) );
  CFD2QXL \Poly7_reg[208]  ( .D(n9896), .CP(clk), .CD(n18332), .Q(
        poly7_shifted[220]) );
  CFD2QXL \Poly7_reg[220]  ( .D(n9884), .CP(clk), .CD(n18332), .Q(
        poly7_shifted[232]) );
  CFD2QXL \Poly7_reg[232]  ( .D(n9872), .CP(clk), .CD(n18332), .Q(
        poly7_shifted[244]) );
  CFD2QXL \Poly7_reg[213]  ( .D(n9891), .CP(clk), .CD(n18332), .Q(
        poly7_shifted[225]) );
  CFD2QXL \Poly7_reg[225]  ( .D(n9879), .CP(clk), .CD(n18333), .Q(
        poly7_shifted[237]) );
  CFD2QXL \Poly7_reg[251]  ( .D(n9853), .CP(clk), .CD(n18333), .Q(
        poly7_shifted[263]) );
  CFD2QXL \Poly7_reg[263]  ( .D(n9841), .CP(clk), .CD(n18333), .Q(
        poly7_shifted[275]) );
  CFD2QXL \Poly7_reg[275]  ( .D(n9829), .CP(clk), .CD(n18333), .Q(
        poly7_shifted[287]) );
  CFD2QXL \Poly7_reg[287]  ( .D(n9817), .CP(clk), .CD(n18333), .Q(
        poly7_shifted[299]) );
  CFD2QXL \Poly7_reg[299]  ( .D(n9805), .CP(clk), .CD(n18333), .Q(
        poly7_shifted[311]) );
  CFD2QXL \Poly7_reg[311]  ( .D(n9793), .CP(clk), .CD(n18333), .Q(
        poly7_shifted[323]) );
  CFD2QXL \Poly7_reg[323]  ( .D(n9781), .CP(clk), .CD(n18333), .Q(
        poly7_shifted[335]) );
  CFD2QXL \Poly7_reg[335]  ( .D(n9769), .CP(clk), .CD(n18333), .Q(
        poly7_shifted[347]) );
  CFD2QXL \Poly7_reg[347]  ( .D(n9757), .CP(clk), .CD(n18333), .Q(
        poly7_shifted[359]) );
  CFD2QXL \Poly7_reg[359]  ( .D(n9745), .CP(clk), .CD(n18333), .Q(
        poly7_shifted[371]) );
  CFD2QXL \Poly7_reg[371]  ( .D(n9733), .CP(clk), .CD(n18333), .Q(
        poly7_shifted[383]) );
  CFD2QXL \Poly7_reg[383]  ( .D(n9721), .CP(clk), .CD(n18333), .Q(
        poly7_shifted[395]) );
  CFD2QXL \Poly7_reg[395]  ( .D(n9709), .CP(clk), .CD(n18333), .Q(
        poly7_shifted[407]) );
  CFD2QXL \Poly7_reg[8]  ( .D(n10096), .CP(clk), .CD(n18334), .Q(
        poly7_shifted[20]) );
  CFD2QXL \Poly7_reg[44]  ( .D(n10060), .CP(clk), .CD(n18334), .Q(
        poly7_shifted[56]) );
  CFD2QXL \Poly7_reg[75]  ( .D(n10029), .CP(clk), .CD(n18334), .Q(
        poly7_shifted[87]) );
  CFD2QXL \Poly7_reg[87]  ( .D(n10017), .CP(clk), .CD(n18334), .Q(
        poly7_shifted[99]) );
  CFD2QXL \Poly7_reg[99]  ( .D(n10005), .CP(clk), .CD(n18334), .Q(
        poly7_shifted[111]) );
  CFD2QXL \Poly7_reg[111]  ( .D(n9993), .CP(clk), .CD(n18334), .Q(
        poly7_shifted[123]) );
  CFD2QXL \Poly7_reg[123]  ( .D(n9981), .CP(clk), .CD(n18334), .Q(
        poly7_shifted[135]) );
  CFD2QXL \Poly7_reg[135]  ( .D(n9969), .CP(clk), .CD(n18334), .Q(
        poly7_shifted[147]) );
  CFD2QXL \Poly7_reg[171]  ( .D(n9933), .CP(clk), .CD(n18334), .Q(
        poly7_shifted[183]) );
  CFD2QXL \Poly7_reg[80]  ( .D(n10024), .CP(clk), .CD(n18335), .Q(
        poly7_shifted[92]) );
  CFD2QXL \Poly7_reg[116]  ( .D(n9988), .CP(clk), .CD(n18335), .Q(
        poly7_shifted[128]) );
  CFD2QXL \Poly7_reg[128]  ( .D(n9976), .CP(clk), .CD(n18335), .Q(
        poly7_shifted[140]) );
  CFD2QXL \Poly7_reg[176]  ( .D(n9928), .CP(clk), .CD(n18335), .Q(
        poly7_shifted[188]) );
  CFD2QXL \Poly7_reg[210]  ( .D(n9894), .CP(clk), .CD(n18335), .Q(
        poly7_shifted[222]) );
  CFD2QXL \Poly7_reg[215]  ( .D(n9889), .CP(clk), .CD(n18336), .Q(
        poly7_shifted[227]) );
  CFD2QXL \Poly7_reg[227]  ( .D(n9877), .CP(clk), .CD(n18336), .Q(
        poly7_shifted[239]) );
  CFD2QXL \Poly7_reg[253]  ( .D(n9851), .CP(clk), .CD(n18336), .Q(
        poly7_shifted[265]) );
  CFD2QXL \Poly7_reg[265]  ( .D(n9839), .CP(clk), .CD(n18336), .Q(
        poly7_shifted[277]) );
  CFD2QXL \Poly7_reg[277]  ( .D(n9827), .CP(clk), .CD(n18336), .Q(
        poly7_shifted[289]) );
  CFD2QXL \Poly7_reg[289]  ( .D(n9815), .CP(clk), .CD(n18336), .Q(
        poly7_shifted[301]) );
  CFD2QXL \Poly7_reg[301]  ( .D(n9803), .CP(clk), .CD(n18336), .Q(
        poly7_shifted[313]) );
  CFD2QXL \Poly7_reg[313]  ( .D(n9791), .CP(clk), .CD(n18336), .Q(
        poly7_shifted[325]) );
  CFD2QXL \Poly7_reg[325]  ( .D(n9779), .CP(clk), .CD(n18336), .Q(
        poly7_shifted[337]) );
  CFD2QXL \Poly7_reg[373]  ( .D(n9731), .CP(clk), .CD(n18336), .Q(
        poly7_shifted[385]) );
  CFD2QXL \Poly7_reg[385]  ( .D(n9719), .CP(clk), .CD(n18336), .Q(
        poly7_shifted[397]) );
  CFD2QXL \Poly7_reg[397]  ( .D(n9707), .CP(clk), .CD(n18336), .Q(
        poly7_shifted[409]) );
  CFD2QXL \Poly7_reg[10]  ( .D(n10094), .CP(clk), .CD(n18337), .Q(
        poly7_shifted[22]) );
  CFD2QXL \Poly7_reg[77]  ( .D(n10027), .CP(clk), .CD(n18337), .Q(
        poly7_shifted[89]) );
  CFD2QXL \Poly7_reg[89]  ( .D(n10015), .CP(clk), .CD(n18337), .Q(
        poly7_shifted[101]) );
  CFD2QXL \Poly7_reg[101]  ( .D(n10003), .CP(clk), .CD(n18337), .Q(
        poly7_shifted[113]) );
  CFD2QXL \Poly7_reg[113]  ( .D(n9991), .CP(clk), .CD(n18337), .Q(
        poly7_shifted[125]) );
  CFD2QXL \Poly7_reg[125]  ( .D(n9979), .CP(clk), .CD(n18337), .Q(
        poly7_shifted[137]) );
  CFD2QXL \Poly7_reg[137]  ( .D(n9967), .CP(clk), .CD(n18337), .Q(
        poly7_shifted[149]) );
  CFD2QXL \Poly7_reg[149]  ( .D(n9955), .CP(clk), .CD(n18337), .Q(
        poly7_shifted[161]) );
  CFD2QXL \Poly7_reg[161]  ( .D(n9943), .CP(clk), .CD(n18337), .Q(
        poly7_shifted[173]) );
  CFD2QXL \Poly7_reg[173]  ( .D(n9931), .CP(clk), .CD(n18337), .Q(
        poly7_shifted[185]) );
  CFD2QXL \Poly7_reg[82]  ( .D(n10022), .CP(clk), .CD(n18338), .Q(
        poly7_shifted[94]) );
  CFD2QXL \Poly7_reg[94]  ( .D(n10010), .CP(clk), .CD(n18338), .Q(
        poly7_shifted[106]) );
  CFD2QXL \Poly7_reg[106]  ( .D(n9998), .CP(clk), .CD(n18338), .Q(
        poly7_shifted[118]) );
  CFD2QXL \Poly7_reg[130]  ( .D(n9974), .CP(clk), .CD(n18338), .Q(
        poly7_shifted[142]) );
  CFD2QXL \Poly7_reg[142]  ( .D(n9962), .CP(clk), .CD(n18338), .Q(
        poly7_shifted[154]) );
  CFD2QXL \Poly7_reg[154]  ( .D(n9950), .CP(clk), .CD(n18338), .Q(
        poly7_shifted[166]) );
  CFD2QXL \Poly7_reg[166]  ( .D(n9938), .CP(clk), .CD(n18338), .Q(
        poly7_shifted[178]) );
  CFD2QXL \Poly7_reg[217]  ( .D(n9887), .CP(clk), .CD(n18338), .Q(
        poly7_shifted[229]) );
  CFD2QXL \Poly7_reg[229]  ( .D(n9875), .CP(clk), .CD(n18339), .Q(
        poly7_shifted[241]) );
  CFD2QXL \Poly7_reg[279]  ( .D(n9825), .CP(clk), .CD(n18339), .Q(
        poly7_shifted[291]) );
  CFD2QXL \Poly7_reg[291]  ( .D(n9813), .CP(clk), .CD(n18339), .Q(
        poly7_shifted[303]) );
  CFD2QXL \Poly7_reg[363]  ( .D(n9741), .CP(clk), .CD(n18339), .Q(
        poly7_shifted[375]) );
  CFD2QXL \Poly7_reg[375]  ( .D(n9729), .CP(clk), .CD(n18339), .Q(
        poly7_shifted[387]) );
  CFD2QXL \Poly7_reg[387]  ( .D(n9717), .CP(clk), .CD(n18339), .Q(
        poly7_shifted[399]) );
  CFD2QXL \Poly7_reg[79]  ( .D(n10025), .CP(clk), .CD(n18340), .Q(
        poly7_shifted[91]) );
  CFD2QXL \Poly7_reg[91]  ( .D(n10013), .CP(clk), .CD(n18340), .Q(
        poly7_shifted[103]) );
  CFD2QXL \Poly7_reg[127]  ( .D(n9977), .CP(clk), .CD(n18340), .Q(
        poly7_shifted[139]) );
  CFD2QXL \Poly7_reg[139]  ( .D(n9965), .CP(clk), .CD(n18340), .Q(
        poly7_shifted[151]) );
  CFD2QXL \Poly7_reg[151]  ( .D(n9953), .CP(clk), .CD(n18340), .Q(
        poly7_shifted[163]) );
  CFD2QXL \Poly7_reg[163]  ( .D(n9941), .CP(clk), .CD(n18340), .Q(
        poly7_shifted[175]) );
  CFD2QXL \Poly7_reg[175]  ( .D(n9929), .CP(clk), .CD(n18340), .Q(
        poly7_shifted[187]) );
  CFD2QXL \Poly7_reg[211]  ( .D(n9893), .CP(clk), .CD(n18340), .Q(
        poly7_shifted[223]) );
  CFD2QXL \Poly7_reg[223]  ( .D(n9881), .CP(clk), .CD(n18340), .Q(
        poly7_shifted[235]) );
  CFD2QXL \Poly7_reg[207]  ( .D(n9897), .CP(clk), .CD(n18341), .Q(
        poly7_shifted[219]) );
  CFD2QXL \Poly7_reg[219]  ( .D(n9885), .CP(clk), .CD(n18341), .Q(
        poly7_shifted[231]) );
  CFD2QXL \Poly7_reg[214]  ( .D(n9890), .CP(clk), .CD(n18341), .Q(
        poly7_shifted[226]) );
  CFD2QXL \Poly7_reg[226]  ( .D(n9878), .CP(clk), .CD(n18341), .Q(
        poly7_shifted[238]) );
  CFD2QXL \Poly15_reg[38]  ( .D(n9599), .CP(clk), .CD(n18345), .Q(
        poly15_shifted[53]) );
  CFD2QXL \Poly15_reg[41]  ( .D(n9596), .CP(clk), .CD(n18346), .Q(
        poly15_shifted[56]) );
  CFD2QXL \Poly15_reg[11]  ( .D(n9626), .CP(clk), .CD(n18346), .Q(
        poly15_shifted[26]) );
  CFD2QXL \Poly15_reg[6]  ( .D(n9631), .CP(clk), .CD(n18256), .Q(
        poly15_shifted[21]) );
  CFD2QXL \Poly1_reg[77]  ( .D(n9280), .CP(clk), .CD(n18358), .Q(
        poly1_shifted[88]) );
  CFD2QXL \Poly1_reg[88]  ( .D(n9269), .CP(clk), .CD(n18358), .Q(
        poly1_shifted[99]) );
  CFD2QXL \Poly1_reg[99]  ( .D(n9258), .CP(clk), .CD(n18358), .Q(
        poly1_shifted[110]) );
  CFD2QXL \Poly1_reg[110]  ( .D(n9247), .CP(clk), .CD(n18358), .Q(
        poly1_shifted[121]) );
  CFD2QXL \Poly1_reg[132]  ( .D(n9225), .CP(clk), .CD(n18359), .Q(
        poly1_shifted[143]) );
  CFD2QXL \Poly1_reg[143]  ( .D(n9214), .CP(clk), .CD(n18359), .Q(
        poly1_shifted[154]) );
  CFD2QXL \Poly1_reg[165]  ( .D(n9192), .CP(clk), .CD(n18359), .Q(
        poly1_shifted[176]) );
  CFD2QXL \Poly1_reg[176]  ( .D(n9181), .CP(clk), .CD(n18359), .Q(
        poly1_shifted[187]) );
  CFD2QXL \Poly1_reg[187]  ( .D(n9170), .CP(clk), .CD(n18359), .Q(
        poly1_shifted[198]) );
  CFD2QXL \Poly1_reg[220]  ( .D(n9137), .CP(clk), .CD(n18359), .Q(
        poly1_shifted[231]) );
  CFD2QXL \Poly1_reg[253]  ( .D(n9104), .CP(clk), .CD(n18359), .Q(
        poly1_shifted[264]) );
  CFD2QXL \Poly1_reg[275]  ( .D(n9082), .CP(clk), .CD(n18359), .Q(
        poly1_shifted[286]) );
  CFD2QXL \Poly1_reg[286]  ( .D(n9071), .CP(clk), .CD(n18359), .Q(
        poly1_shifted[297]) );
  CFD2QXL \Poly1_reg[297]  ( .D(n9060), .CP(clk), .CD(n18359), .Q(
        poly1_shifted[308]) );
  CFD2QXL \Poly1_reg[330]  ( .D(n9027), .CP(clk), .CD(n18360), .Q(
        poly1_shifted[341]) );
  CFD2QXL \Poly1_reg[263]  ( .D(n9094), .CP(clk), .CD(n18360), .Q(
        poly1_shifted[274]) );
  CFD2QXL \Poly1_reg[274]  ( .D(n9083), .CP(clk), .CD(n18360), .Q(
        poly1_shifted[285]) );
  CFD2QXL \Poly1_reg[296]  ( .D(n9061), .CP(clk), .CD(n18360), .Q(
        poly1_shifted[307]) );
  CFD2QXL \Poly1_reg[318]  ( .D(n9039), .CP(clk), .CD(n18360), .Q(
        poly1_shifted[329]) );
  CFD2QXL \Poly1_reg[329]  ( .D(n9028), .CP(clk), .CD(n18360), .Q(
        poly1_shifted[340]) );
  CFD2QXL \Poly1_reg[251]  ( .D(n9106), .CP(clk), .CD(n18361), .Q(
        poly1_shifted[262]) );
  CFD2QXL \Poly1_reg[262]  ( .D(n9095), .CP(clk), .CD(n18361), .Q(
        poly1_shifted[273]) );
  CFD2QXL \Poly1_reg[273]  ( .D(n9084), .CP(clk), .CD(n18361), .Q(
        poly1_shifted[284]) );
  CFD2QXL \Poly1_reg[306]  ( .D(n9051), .CP(clk), .CD(n18361), .Q(
        poly1_shifted[317]) );
  CFD2QXL \Poly1_reg[317]  ( .D(n9040), .CP(clk), .CD(n18361), .Q(
        poly1_shifted[328]) );
  CFD2QXL \Poly1_reg[328]  ( .D(n9029), .CP(clk), .CD(n18361), .Q(
        poly1_shifted[339]) );
  CFD2QXL \Poly1_reg[80]  ( .D(n9277), .CP(clk), .CD(n18362), .Q(
        poly1_shifted[91]) );
  CFD2QXL \Poly1_reg[91]  ( .D(n9266), .CP(clk), .CD(n18362), .Q(
        poly1_shifted[102]) );
  CFD2QXL \Poly1_reg[102]  ( .D(n9255), .CP(clk), .CD(n18362), .Q(
        poly1_shifted[113]) );
  CFD2QXL \Poly1_reg[113]  ( .D(n9244), .CP(clk), .CD(n18362), .Q(
        poly1_shifted[124]) );
  CFD2QXL \Poly1_reg[124]  ( .D(n9233), .CP(clk), .CD(n18362), .Q(
        poly1_shifted[135]) );
  CFD2QXL \Poly1_reg[135]  ( .D(n9222), .CP(clk), .CD(n18362), .Q(
        poly1_shifted[146]) );
  CFD2QXL \Poly1_reg[146]  ( .D(n9211), .CP(clk), .CD(n18362), .Q(
        poly1_shifted[157]) );
  CFD2QXL \Poly1_reg[239]  ( .D(n9118), .CP(clk), .CD(n18362), .Q(
        poly1_shifted[250]) );
  CFD2QXL \Poly1_reg[250]  ( .D(n9107), .CP(clk), .CD(n18362), .Q(
        poly1_shifted[261]) );
  CFD2QXL \Poly1_reg[261]  ( .D(n9096), .CP(clk), .CD(n18362), .Q(
        poly1_shifted[272]) );
  CFD2QXL \Poly1_reg[272]  ( .D(n9085), .CP(clk), .CD(n18362), .Q(
        poly1_shifted[283]) );
  CFD2QXL \Poly1_reg[283]  ( .D(n9074), .CP(clk), .CD(n18362), .Q(
        poly1_shifted[294]) );
  CFD2QXL \Poly1_reg[316]  ( .D(n9041), .CP(clk), .CD(n18363), .Q(
        poly1_shifted[327]) );
  CFD2QXL \Poly1_reg[327]  ( .D(n9030), .CP(clk), .CD(n18363), .Q(
        poly1_shifted[338]) );
  CFD2QXL \Poly1_reg[46]  ( .D(n9311), .CP(clk), .CD(n18363), .Q(
        poly1_shifted[57]) );
  CFD2QXL \Poly1_reg[79]  ( .D(n9278), .CP(clk), .CD(n18363), .Q(
        poly1_shifted[90]) );
  CFD2QXL \Poly1_reg[101]  ( .D(n9256), .CP(clk), .CD(n18363), .Q(
        poly1_shifted[112]) );
  CFD2QXL \Poly1_reg[112]  ( .D(n9245), .CP(clk), .CD(n18363), .Q(
        poly1_shifted[123]) );
  CFD2QXL \Poly1_reg[123]  ( .D(n9234), .CP(clk), .CD(n18363), .Q(
        poly1_shifted[134]) );
  CFD2QXL \Poly1_reg[260]  ( .D(n9097), .CP(clk), .CD(n18364), .Q(
        poly1_shifted[271]) );
  CFD2QXL \Poly1_reg[271]  ( .D(n9086), .CP(clk), .CD(n18364), .Q(
        poly1_shifted[282]) );
  CFD2QXL \Poly1_reg[282]  ( .D(n9075), .CP(clk), .CD(n18364), .Q(
        poly1_shifted[293]) );
  CFD2QXL \Poly1_reg[293]  ( .D(n9064), .CP(clk), .CD(n18364), .Q(
        poly1_shifted[304]) );
  CFD2QXL \Poly1_reg[315]  ( .D(n9042), .CP(clk), .CD(n18364), .Q(
        poly1_shifted[326]) );
  CFD2QXL \Poly1_reg[326]  ( .D(n9031), .CP(clk), .CD(n18364), .Q(
        poly1_shifted[337]) );
  CFD2QXL \Poly1_reg[34]  ( .D(n9323), .CP(clk), .CD(n18365), .Q(
        poly1_shifted[45]) );
  CFD2QXL \Poly1_reg[45]  ( .D(n9312), .CP(clk), .CD(n18365), .Q(
        poly1_shifted[56]) );
  CFD2QXL \Poly1_reg[67]  ( .D(n9290), .CP(clk), .CD(n18365), .Q(
        poly1_shifted[78]) );
  CFD2QXL \Poly1_reg[78]  ( .D(n9279), .CP(clk), .CD(n18365), .Q(
        poly1_shifted[89]) );
  CFD2QXL \Poly1_reg[100]  ( .D(n9257), .CP(clk), .CD(n18365), .Q(
        poly1_shifted[111]) );
  CFD2QXL \Poly1_reg[111]  ( .D(n9246), .CP(clk), .CD(n18365), .Q(
        poly1_shifted[122]) );
  CFD2QXL \Poly1_reg[122]  ( .D(n9235), .CP(clk), .CD(n18365), .Q(
        poly1_shifted[133]) );
  CFD2QXL \Poly1_reg[133]  ( .D(n9224), .CP(clk), .CD(n18365), .Q(
        poly1_shifted[144]) );
  CFD2QXL \Poly1_reg[144]  ( .D(n9213), .CP(clk), .CD(n18365), .Q(
        poly1_shifted[155]) );
  CFD2QXL \Poly1_reg[188]  ( .D(n9169), .CP(clk), .CD(n18365), .Q(
        poly1_shifted[199]) );
  CFD2QXL \Poly1_reg[221]  ( .D(n9136), .CP(clk), .CD(n18254), .Q(
        poly1_shifted[232]) );
  CFD2QXL \Poly1_reg[259]  ( .D(n9098), .CP(clk), .CD(n18254), .Q(
        poly1_shifted[270]) );
  CFD2QXL \Poly1_reg[270]  ( .D(n9087), .CP(clk), .CD(n18254), .Q(
        poly1_shifted[281]) );
  CFD2QXL \Poly1_reg[281]  ( .D(n9076), .CP(clk), .CD(n18254), .Q(
        poly1_shifted[292]) );
  CFD2QXL \Poly1_reg[292]  ( .D(n9065), .CP(clk), .CD(n18254), .Q(
        poly1_shifted[303]) );
  CFD2QXL \Poly1_reg[303]  ( .D(n9054), .CP(clk), .CD(n18254), .Q(
        poly1_shifted[314]) );
  CFD2QXL \Poly1_reg[314]  ( .D(n9043), .CP(clk), .CD(n18254), .Q(
        poly1_shifted[325]) );
  CFD2QXL \Poly1_reg[325]  ( .D(n9032), .CP(clk), .CD(n18254), .Q(
        poly1_shifted[336]) );
  CFD2QXL \Poly1_reg[258]  ( .D(n9099), .CP(clk), .CD(n18254), .Q(
        poly1_shifted[269]) );
  CFD2QXL \Poly1_reg[269]  ( .D(n9088), .CP(clk), .CD(n18366), .Q(
        poly1_shifted[280]) );
  CFD2QXL \Poly1_reg[280]  ( .D(n9077), .CP(clk), .CD(n18366), .Q(
        poly1_shifted[291]) );
  CFD2QXL \Poly1_reg[291]  ( .D(n9066), .CP(clk), .CD(n18366), .Q(
        poly1_shifted[302]) );
  CFD2QXL \Poly1_reg[324]  ( .D(n9033), .CP(clk), .CD(n18366), .Q(
        poly1_shifted[335]) );
  CFD2QXL \Poly1_reg[335]  ( .D(n9022), .CP(clk), .CD(n18366), .Q(
        poly1_shifted[346]) );
  CFD2QXL \Poly1_reg[43]  ( .D(n9314), .CP(clk), .CD(n18366), .Q(
        poly1_shifted[54]) );
  CFD2QXL \Poly1_reg[76]  ( .D(n9281), .CP(clk), .CD(n18366), .Q(
        poly1_shifted[87]) );
  CFD2QXL \Poly1_reg[87]  ( .D(n9270), .CP(clk), .CD(n18366), .Q(
        poly1_shifted[98]) );
  CFD2QXL \Poly1_reg[98]  ( .D(n9259), .CP(clk), .CD(n18366), .Q(
        poly1_shifted[109]) );
  CFD2QXL \Poly1_reg[109]  ( .D(n9248), .CP(clk), .CD(n18366), .Q(
        poly1_shifted[120]) );
  CFD2QXL \Poly1_reg[142]  ( .D(n9215), .CP(clk), .CD(n18367), .Q(
        poly1_shifted[153]) );
  CFD2QXL \Poly1_reg[175]  ( .D(n9182), .CP(clk), .CD(n18367), .Q(
        poly1_shifted[186]) );
  CFD2QXL \Poly1_reg[186]  ( .D(n9171), .CP(clk), .CD(n18367), .Q(
        poly1_shifted[197]) );
  CFD2QXL \Poly1_reg[197]  ( .D(n9160), .CP(clk), .CD(n18367), .Q(
        poly1_shifted[208]) );
  CFD2QXL \Poly1_reg[219]  ( .D(n9138), .CP(clk), .CD(n18367), .Q(
        poly1_shifted[230]) );
  CFD2QXL \Poly1_reg[257]  ( .D(n9100), .CP(clk), .CD(n18367), .Q(
        poly1_shifted[268]) );
  CFD2QXL \Poly1_reg[268]  ( .D(n9089), .CP(clk), .CD(n18367), .Q(
        poly1_shifted[279]) );
  CFD2QXL \Poly1_reg[301]  ( .D(n9056), .CP(clk), .CD(n18367), .Q(
        poly1_shifted[312]) );
  CFD2QXL \Poly1_reg[312]  ( .D(n9045), .CP(clk), .CD(n18368), .Q(
        poly1_shifted[323]) );
  CFD2QXL \Poly1_reg[323]  ( .D(n9034), .CP(clk), .CD(n18368), .Q(
        poly1_shifted[334]) );
  CFD2QXL \Poly1_reg[334]  ( .D(n9023), .CP(clk), .CD(n18368), .Q(
        poly1_shifted[345]) );
  CFD2QXL \Poly1_reg[75]  ( .D(n9282), .CP(clk), .CD(n18368), .Q(
        poly1_shifted[86]) );
  CFD2QXL \Poly1_reg[86]  ( .D(n9271), .CP(clk), .CD(n18368), .Q(
        poly1_shifted[97]) );
  CFD2QXL \Poly1_reg[97]  ( .D(n9260), .CP(clk), .CD(n18368), .Q(
        poly1_shifted[108]) );
  CFD2QXL \Poly1_reg[108]  ( .D(n9249), .CP(clk), .CD(n18368), .Q(
        poly1_shifted[119]) );
  CFD2QXL \Poly1_reg[119]  ( .D(n9238), .CP(clk), .CD(n18368), .Q(
        poly1_shifted[130]) );
  CFD2QXL \Poly1_reg[130]  ( .D(n9227), .CP(clk), .CD(n18368), .Q(
        poly1_shifted[141]) );
  CFD2QXL \Poly1_reg[141]  ( .D(n9216), .CP(clk), .CD(n18368), .Q(
        poly1_shifted[152]) );
  CFD2QXL \Poly1_reg[185]  ( .D(n9172), .CP(clk), .CD(n18369), .Q(
        poly1_shifted[196]) );
  CFD2QXL \Poly1_reg[196]  ( .D(n9161), .CP(clk), .CD(n18369), .Q(
        poly1_shifted[207]) );
  CFD2QXL \Poly1_reg[278]  ( .D(n9079), .CP(clk), .CD(n18369), .Q(
        poly1_shifted[289]) );
  CFD2QXL \Poly1_reg[311]  ( .D(n9046), .CP(clk), .CD(n18369), .Q(
        poly1_shifted[322]) );
  CFD2QXL \Poly1_reg[322]  ( .D(n9035), .CP(clk), .CD(n18369), .Q(
        poly1_shifted[333]) );
  CFD2QXL \Poly1_reg[333]  ( .D(n9024), .CP(clk), .CD(n18370), .Q(
        poly1_shifted[344]) );
  CFD2QXL \Poly1_reg[52]  ( .D(n9305), .CP(clk), .CD(n18370), .Q(
        poly1_shifted[63]) );
  CFD2QXL \Poly1_reg[107]  ( .D(n9250), .CP(clk), .CD(n18370), .Q(
        poly1_shifted[118]) );
  CFD2QXL \Poly1_reg[118]  ( .D(n9239), .CP(clk), .CD(n18370), .Q(
        poly1_shifted[129]) );
  CFD2QXL \Poly1_reg[129]  ( .D(n9228), .CP(clk), .CD(n18370), .Q(
        poly1_shifted[140]) );
  CFD2QXL \Poly1_reg[140]  ( .D(n9217), .CP(clk), .CD(n18370), .Q(
        poly1_shifted[151]) );
  CFD2QXL \Poly1_reg[184]  ( .D(n9173), .CP(clk), .CD(n18371), .Q(
        poly1_shifted[195]) );
  CFD2QXL \Poly1_reg[195]  ( .D(n9162), .CP(clk), .CD(n18371), .Q(
        poly1_shifted[206]) );
  CFD2QXL \Poly1_reg[266]  ( .D(n9091), .CP(clk), .CD(n18371), .Q(
        poly1_shifted[277]) );
  CFD2QXL \Poly1_reg[277]  ( .D(n9080), .CP(clk), .CD(n18371), .Q(
        poly1_shifted[288]) );
  CFD2QXL \Poly1_reg[299]  ( .D(n9058), .CP(clk), .CD(n18371), .Q(
        poly1_shifted[310]) );
  CFD2QXL \Poly1_reg[310]  ( .D(n9047), .CP(clk), .CD(n18371), .Q(
        poly1_shifted[321]) );
  CFD2QXL \Poly1_reg[321]  ( .D(n9036), .CP(clk), .CD(n18371), .Q(
        poly1_shifted[332]) );
  CFD2QXL \Poly1_reg[332]  ( .D(n9025), .CP(clk), .CD(n18371), .Q(
        poly1_shifted[343]) );
  CFD2QXL \Poly1_reg[51]  ( .D(n9306), .CP(clk), .CD(n18372), .Q(
        poly1_shifted[62]) );
  CFD2QXL \Poly1_reg[84]  ( .D(n9273), .CP(clk), .CD(n18372), .Q(
        poly1_shifted[95]) );
  CFD2QXL \Poly1_reg[95]  ( .D(n9262), .CP(clk), .CD(n18372), .Q(
        poly1_shifted[106]) );
  CFD2QXL \Poly1_reg[106]  ( .D(n9251), .CP(clk), .CD(n18372), .Q(
        poly1_shifted[117]) );
  CFD2QXL \Poly1_reg[117]  ( .D(n9240), .CP(clk), .CD(n18372), .Q(
        poly1_shifted[128]) );
  CFD2QXL \Poly1_reg[128]  ( .D(n9229), .CP(clk), .CD(n18372), .Q(
        poly1_shifted[139]) );
  CFD2QXL \Poly1_reg[139]  ( .D(n9218), .CP(clk), .CD(n18372), .Q(
        poly1_shifted[150]) );
  CFD2QXL \Poly1_reg[150]  ( .D(n9207), .CP(clk), .CD(n18372), .Q(
        poly1_shifted[161]) );
  CFD2QXL \Poly1_reg[183]  ( .D(n9174), .CP(clk), .CD(n18372), .Q(
        poly1_shifted[194]) );
  CFD2QXL \Poly1_reg[194]  ( .D(n9163), .CP(clk), .CD(n18372), .Q(
        poly1_shifted[205]) );
  CFD2QXL \Poly1_reg[82]  ( .D(n9275), .CP(clk), .CD(n18373), .Q(
        poly1_shifted[93]) );
  CFD2QXL \Poly1_reg[93]  ( .D(n9264), .CP(clk), .CD(n18373), .Q(
        poly1_shifted[104]) );
  CFD2QXL \Poly1_reg[104]  ( .D(n9253), .CP(clk), .CD(n18373), .Q(
        poly1_shifted[115]) );
  CFD2QXL \Poly1_reg[115]  ( .D(n9242), .CP(clk), .CD(n18373), .Q(
        poly1_shifted[126]) );
  CFD2QXL \Poly1_reg[126]  ( .D(n9231), .CP(clk), .CD(n18373), .Q(
        poly1_shifted[137]) );
  CFD2QXL \Poly1_reg[137]  ( .D(n9220), .CP(clk), .CD(n18373), .Q(
        poly1_shifted[148]) );
  CFD2QXL \Poly1_reg[148]  ( .D(n9209), .CP(clk), .CD(n18373), .Q(
        poly1_shifted[159]) );
  CFD2QXL \Poly1_reg[181]  ( .D(n9176), .CP(clk), .CD(n18373), .Q(
        poly1_shifted[192]) );
  CFD2QXL \Poly1_reg[192]  ( .D(n9165), .CP(clk), .CD(n18373), .Q(
        poly1_shifted[203]) );
  CFD2QXL \Poly1_reg[276]  ( .D(n9081), .CP(clk), .CD(n18374), .Q(
        poly1_shifted[287]) );
  CFD2QXL \Poly1_reg[287]  ( .D(n9070), .CP(clk), .CD(n18374), .Q(
        poly1_shifted[298]) );
  CFD2QXL \Poly1_reg[298]  ( .D(n9059), .CP(clk), .CD(n18374), .Q(
        poly1_shifted[309]) );
  CFD2QXL \Poly1_reg[309]  ( .D(n9048), .CP(clk), .CD(n18374), .Q(
        poly1_shifted[320]) );
  CFD2QXL \Poly1_reg[320]  ( .D(n9037), .CP(clk), .CD(n18374), .Q(
        poly1_shifted[331]) );
  CFD2QXL \Poly1_reg[331]  ( .D(n9026), .CP(clk), .CD(n18374), .Q(
        poly1_shifted[342]) );
  CFD2QXL \Poly1_reg[50]  ( .D(n9307), .CP(clk), .CD(n18375), .Q(
        poly1_shifted[61]) );
  CFD2QXL \Poly1_reg[83]  ( .D(n9274), .CP(clk), .CD(n18375), .Q(
        poly1_shifted[94]) );
  CFD2QXL \Poly1_reg[94]  ( .D(n9263), .CP(clk), .CD(n18375), .Q(
        poly1_shifted[105]) );
  CFD2QXL \Poly1_reg[105]  ( .D(n9252), .CP(clk), .CD(n18375), .Q(
        poly1_shifted[116]) );
  CFD2QXL \Poly1_reg[138]  ( .D(n9219), .CP(clk), .CD(n18375), .Q(
        poly1_shifted[149]) );
  CFD2QXL \Poly1_reg[182]  ( .D(n9175), .CP(clk), .CD(n18375), .Q(
        poly1_shifted[193]) );
  CFD2QXL \Poly1_reg[193]  ( .D(n9164), .CP(clk), .CD(n18375), .Q(
        poly1_shifted[204]) );
  CFD2QXL \Poly1_reg[48]  ( .D(n9309), .CP(clk), .CD(n18375), .Q(
        poly1_shifted[59]) );
  CFD2QXL \Poly1_reg[92]  ( .D(n9265), .CP(clk), .CD(n18376), .Q(
        poly1_shifted[103]) );
  CFD2QXL \Poly1_reg[114]  ( .D(n9243), .CP(clk), .CD(n18376), .Q(
        poly1_shifted[125]) );
  CFD2QXL \Poly1_reg[125]  ( .D(n9232), .CP(clk), .CD(n18376), .Q(
        poly1_shifted[136]) );
  CFD2QXL \Poly1_reg[136]  ( .D(n9221), .CP(clk), .CD(n18376), .Q(
        poly1_shifted[147]) );
  CFD2QXL \Poly1_reg[147]  ( .D(n9210), .CP(clk), .CD(n18376), .Q(
        poly1_shifted[158]) );
  CFD2QXL \Poly1_reg[180]  ( .D(n9177), .CP(clk), .CD(n18376), .Q(
        poly1_shifted[191]) );
  CFD2QXL \Poly1_reg[191]  ( .D(n9166), .CP(clk), .CD(n18376), .Q(
        poly1_shifted[202]) );
  CFD2QXL \Poly1_reg[224]  ( .D(n9133), .CP(clk), .CD(n18376), .Q(
        poly1_shifted[235]) );
  CFD2QXL \Poly1_reg[179]  ( .D(n9178), .CP(clk), .CD(n18377), .Q(
        poly1_shifted[190]) );
  CFD2QXL \Poly1_reg[190]  ( .D(n9167), .CP(clk), .CD(n18377), .Q(
        poly1_shifted[201]) );
  CFD2QXL \Poly1_reg[212]  ( .D(n9145), .CP(clk), .CD(n18377), .Q(
        poly1_shifted[223]) );
  CFD2QXL \Poly1_reg[223]  ( .D(n9134), .CP(clk), .CD(n18377), .Q(
        poly1_shifted[234]) );
  CFD2QXL \Poly2_reg[0]  ( .D(n9010), .CP(clk), .CD(n18377), .Q(
        poly2_shifted[12]) );
  CFD2QXL \Poly2_reg[12]  ( .D(n8998), .CP(clk), .CD(n18377), .Q(
        poly2_shifted[24]) );
  CFD2QXL \Poly2_reg[2]  ( .D(n9008), .CP(clk), .CD(n18377), .Q(
        poly2_shifted[14]) );
  CFD2QXL \Poly2_reg[14]  ( .D(n8996), .CP(clk), .CD(n18377), .Q(
        poly2_shifted[26]) );
  CFD2QXL \Poly2_reg[9]  ( .D(n9001), .CP(clk), .CD(n18378), .Q(
        poly2_shifted[21]) );
  CFD2QXL \Poly2_reg[6]  ( .D(n9004), .CP(clk), .CD(n18378), .Q(
        poly2_shifted[18]) );
  CFD2QXL \Poly2_reg[10]  ( .D(n9000), .CP(clk), .CD(n18379), .Q(
        poly2_shifted[22]) );
  CFD2QXL \Poly2_reg[15]  ( .D(n8995), .CP(clk), .CD(n18379), .Q(
        poly2_shifted[27]) );
  CFD2QXL \Poly3_reg[0]  ( .D(n8940), .CP(clk), .CD(n18380), .Q(
        poly3_shifted[14]) );
  CFD2QXL \Poly3_reg[14]  ( .D(n8926), .CP(clk), .CD(n18380), .Q(
        poly3_shifted[28]) );
  CFD2QXL \Poly3_reg[17]  ( .D(n8923), .CP(clk), .CD(n18380), .Q(
        poly3_shifted[31]) );
  CFD2QXL \Poly3_reg[26]  ( .D(n8914), .CP(clk), .CD(n18381), .Q(
        poly3_shifted[40]) );
  CFD2QXL \Poly3_reg[29]  ( .D(n8911), .CP(clk), .CD(n18382), .Q(
        poly3_shifted[43]) );
  CFD2QXL \Poly3_reg[4]  ( .D(n8936), .CP(clk), .CD(n18382), .Q(
        poly3_shifted[18]) );
  CFD2QXL \Poly3_reg[18]  ( .D(n8922), .CP(clk), .CD(n18382), .Q(
        poly3_shifted[32]) );
  CFD2QXL \Poly3_reg[21]  ( .D(n8919), .CP(clk), .CD(n18382), .Q(
        poly3_shifted[35]) );
  CFD2QXL \Poly3_reg[10]  ( .D(n8930), .CP(clk), .CD(n18383), .Q(
        poly3_shifted[24]) );
  CFD2QXL \Poly3_reg[24]  ( .D(n8916), .CP(clk), .CD(n18383), .Q(
        poly3_shifted[38]) );
  CFD2QXL \Poly3_reg[2]  ( .D(n8938), .CP(clk), .CD(n18383), .Q(
        poly3_shifted[16]) );
  CFD2QXL \Poly3_reg[16]  ( .D(n8924), .CP(clk), .CD(n18383), .Q(
        poly3_shifted[30]) );
  CFD2QXL \Poly3_reg[5]  ( .D(n8935), .CP(clk), .CD(n18383), .Q(
        poly3_shifted[19]) );
  CFD2QXL \Poly3_reg[19]  ( .D(n8921), .CP(clk), .CD(n18383), .Q(
        poly3_shifted[33]) );
  CFD2QXL \Poly4_reg[13]  ( .D(n8843), .CP(clk), .CD(n18256), .Q(
        poly4_shifted[30]) );
  CFD2QXL \Poly12_reg[15]  ( .D(n10517), .CP(clk), .CD(n18294), .Q(Poly12[15])
         );
  CFD2QXL \Poly12_reg[92]  ( .D(n10440), .CP(clk), .CD(n18296), .Q(Poly12[92])
         );
  CFD2QXL \Poly12_reg[82]  ( .D(n10450), .CP(clk), .CD(n18398), .Q(Poly12[82])
         );
  CFD2QXL \Poly12_reg[85]  ( .D(n10447), .CP(clk), .CD(n18299), .Q(Poly12[85])
         );
  CFD2QXL \Poly7_reg[55]  ( .D(n10049), .CP(clk), .CD(n18340), .Q(Poly7[55])
         );
  CFD2QXL \Poly0_reg[162]  ( .D(n9415), .CP(clk), .CD(n18347), .Q(Poly0[162])
         );
  CFD2QXL \Poly0_reg[164]  ( .D(n9413), .CP(clk), .CD(n18355), .Q(Poly0[164])
         );
  CFD2QXL \Poly0_reg[163]  ( .D(n9414), .CP(clk), .CD(n18357), .Q(Poly0[163])
         );
  CFD2QXL \Poly1_reg[55]  ( .D(n9302), .CP(clk), .CD(n18358), .Q(Poly1[55]) );
  CFD2QXL \Poly2_reg[40]  ( .D(n8970), .CP(clk), .CD(n18391), .Q(Poly2[40]) );
  CFD2QXL \Poly3_reg[51]  ( .D(n8889), .CP(clk), .CD(n18390), .Q(Poly3[51]) );
  CFD2QXL \Poly3_reg[55]  ( .D(n8885), .CP(clk), .CD(n18390), .Q(Poly3[55]) );
  CFD2QXL \Poly0_reg[100]  ( .D(n9477), .CP(clk), .CD(n18351), .Q(
        poly0_shifted[118]) );
  CFD2QXL \Poly0_reg[133]  ( .D(n9444), .CP(clk), .CD(n18349), .Q(
        poly0_shifted[151]) );
  CFD2QXL \Poly0_reg[28]  ( .D(n9549), .CP(clk), .CD(n18351), .Q(
        poly0_shifted[46]) );
  CFD2QXL \Poly0_reg[25]  ( .D(n9552), .CP(clk), .CD(n18351), .Q(
        poly0_shifted[43]) );
  CFD2QXL \Poly0_reg[134]  ( .D(n9443), .CP(clk), .CD(n18354), .Q(
        poly0_shifted[152]) );
  CFD2QXL \Poly0_reg[132]  ( .D(n9445), .CP(clk), .CD(n18358), .Q(
        poly0_shifted[150]) );
  CFD2QXL \Poly3_reg[68]  ( .D(n8872), .CP(clk), .CD(n18381), .Q(
        poly3_shifted[82]) );
  CFD2QXL \Poly5_reg[7]  ( .D(n11519), .CP(clk), .CD(n18259), .Q(
        poly5_shifted[21]) );
  CFD2QXL \polydata_reg[15]  ( .D(n8699), .CP(clk), .CD(n18401), .Q(
        polydata[15]) );
  CFD2QXL \Poly5_reg[42]  ( .D(n11484), .CP(clk), .CD(n18257), .Q(
        poly5_shifted[56]) );
  CFD2QXL \Poly5_reg[30]  ( .D(n11496), .CP(clk), .CD(n18258), .Q(
        poly5_shifted[44]) );
  CFD2QXL \Poly5_reg[58]  ( .D(n11468), .CP(clk), .CD(n18258), .Q(
        poly5_shifted[72]) );
  CFD2QXL \Poly5_reg[21]  ( .D(n11505), .CP(clk), .CD(n18259), .Q(
        poly5_shifted[35]) );
  CFD2QXL \Poly5_reg[50]  ( .D(n11476), .CP(clk), .CD(n18259), .Q(
        poly5_shifted[64]) );
  CFD2QXL \Poly5_reg[55]  ( .D(n11471), .CP(clk), .CD(n18259), .Q(
        poly5_shifted[69]) );
  CFD2QXL \Poly5_reg[61]  ( .D(n11465), .CP(clk), .CD(n18257), .Q(
        poly5_shifted[75]) );
  CFD2QXL \Poly5_reg[53]  ( .D(n11473), .CP(clk), .CD(n18257), .Q(
        poly5_shifted[67]) );
  CFD2QXL \Poly5_reg[73]  ( .D(n11453), .CP(clk), .CD(n18257), .Q(
        poly5_shifted[87]) );
  CFD2QXL \Poly5_reg[23]  ( .D(n11503), .CP(clk), .CD(n18257), .Q(
        poly5_shifted[37]) );
  CFD2QXL \Poly5_reg[51]  ( .D(n11475), .CP(clk), .CD(n18260), .Q(
        poly5_shifted[65]) );
  CFD2QXL \Poly5_reg[29]  ( .D(n11497), .CP(clk), .CD(n18260), .Q(
        poly5_shifted[43]) );
  CFD2QXL \Poly8_reg[81]  ( .D(n11320), .CP(clk), .CD(n18257), .Q(
        poly8_shifted[95]) );
  CFD2QXL \Poly8_reg[31]  ( .D(n11370), .CP(clk), .CD(n18257), .Q(
        poly8_shifted[45]) );
  CFD2QXL \Poly9_reg[7]  ( .D(n11298), .CP(clk), .CD(n18257), .Q(
        poly9_shifted[18]) );
  CFD2QXL \Poly9_reg[8]  ( .D(n11297), .CP(clk), .CD(n18257), .Q(
        poly9_shifted[19]) );
  CFD2QXL \Poly9_reg[67]  ( .D(n11238), .CP(clk), .CD(n18257), .Q(
        poly9_shifted[78]) );
  CFD2QXL \Poly9_reg[79]  ( .D(n11226), .CP(clk), .CD(n18257), .Q(
        poly9_shifted[90]) );
  CFD2QXL \Poly9_reg[52]  ( .D(n11253), .CP(clk), .CD(n18257), .Q(
        poly9_shifted[63]) );
  CFD2QXL \Poly9_reg[53]  ( .D(n11252), .CP(clk), .CD(n18257), .Q(
        poly9_shifted[64]) );
  CFD2QXL \Poly11_reg[4]  ( .D(n11185), .CP(clk), .CD(n18257), .Q(
        poly11_shifted[19]) );
  CFD2QXL \Poly11_reg[8]  ( .D(n11181), .CP(clk), .CD(n18257), .Q(
        poly11_shifted[23]) );
  CFD2QXL \Poly11_reg[7]  ( .D(n11182), .CP(clk), .CD(n18257), .Q(
        poly11_shifted[22]) );
  CFD2QXL \Poly13_reg[154]  ( .D(n10906), .CP(clk), .CD(n18264), .Q(
        poly13_shifted[168]) );
  CFD2QXL \Poly13_reg[432]  ( .D(n10628), .CP(clk), .CD(n18269), .Q(
        poly13_shifted[446]) );
  CFD2QXL \Poly13_reg[255]  ( .D(n10805), .CP(clk), .CD(n18257), .Q(
        poly13_shifted[269]) );
  CFD2QXL \Poly13_reg[127]  ( .D(n10933), .CP(clk), .CD(n18270), .Q(
        poly13_shifted[141]) );
  CFD2QXL \Poly13_reg[352]  ( .D(n10708), .CP(clk), .CD(n18275), .Q(
        poly13_shifted[366]) );
  CFD2QXL \Poly13_reg[110]  ( .D(n10950), .CP(clk), .CD(n18276), .Q(
        poly13_shifted[124]) );
  CFD2QXL \Poly13_reg[365]  ( .D(n10695), .CP(clk), .CD(n18255), .Q(
        poly13_shifted[379]) );
  CFD2QXL \Poly13_reg[425]  ( .D(n10635), .CP(clk), .CD(n18280), .Q(
        poly13_shifted[439]) );
  CFD2QXL \Poly13_reg[495]  ( .D(n10565), .CP(clk), .CD(n18281), .Q(
        poly13_shifted[509]) );
  CFD2QXL \Poly13_reg[133]  ( .D(n10927), .CP(clk), .CD(n18285), .Q(
        poly13_shifted[147]) );
  CFD2QXL \Poly13_reg[450]  ( .D(n10610), .CP(clk), .CD(n18286), .Q(
        poly13_shifted[464]) );
  CFD2QXL \Poly13_reg[313]  ( .D(n10747), .CP(clk), .CD(n18290), .Q(
        poly13_shifted[327]) );
  CFD2QXL \Poly12_reg[5]  ( .D(n10527), .CP(clk), .CD(n18293), .Q(
        poly12_shifted[21]) );
  CFD2QXL \Poly12_reg[13]  ( .D(n10519), .CP(clk), .CD(n18294), .Q(
        poly12_shifted[29]) );
  CFD2QXL \Poly12_reg[47]  ( .D(n10485), .CP(clk), .CD(n18297), .Q(
        poly12_shifted[63]) );
  CFD2QXL \Poly14_reg[51]  ( .D(n10354), .CP(clk), .CD(n18300), .Q(
        poly14_shifted[67]) );
  CFD2QXL \Poly14_reg[234]  ( .D(n10171), .CP(clk), .CD(n18300), .Q(
        poly14_shifted[250]) );
  CFD2QXL \Poly14_reg[65]  ( .D(n10340), .CP(clk), .CD(n18303), .Q(
        poly14_shifted[81]) );
  CFD2QXL \Poly14_reg[242]  ( .D(n10163), .CP(clk), .CD(n18304), .Q(
        poly14_shifted[258]) );
  CFD2QXL \Poly14_reg[73]  ( .D(n10332), .CP(clk), .CD(n18307), .Q(
        poly14_shifted[89]) );
  CFD2QXL \Poly14_reg[118]  ( .D(n10287), .CP(clk), .CD(n18309), .Q(
        poly14_shifted[134]) );
  CFD2QXL \Poly14_reg[78]  ( .D(n10327), .CP(clk), .CD(n18313), .Q(
        poly14_shifted[94]) );
  CFD2QXL \Poly7_reg[290]  ( .D(n9814), .CP(clk), .CD(n18319), .Q(
        poly7_shifted[302]) );
  CFD2QXL \Poly7_reg[330]  ( .D(n9774), .CP(clk), .CD(n18321), .Q(
        poly7_shifted[342]) );
  CFD2QXL \Poly7_reg[390]  ( .D(n9714), .CP(clk), .CD(n18321), .Q(
        poly7_shifted[402]) );
  CFD2QXL \Poly7_reg[158]  ( .D(n9946), .CP(clk), .CD(n18326), .Q(
        poly7_shifted[170]) );
  CFD2QXL \Poly7_reg[379]  ( .D(n9725), .CP(clk), .CD(n18327), .Q(
        poly7_shifted[391]) );
  CFD2QXL \Poly7_reg[230]  ( .D(n9874), .CP(clk), .CD(n18329), .Q(
        poly7_shifted[242]) );
  CFD2QXL \Poly7_reg[85]  ( .D(n10019), .CP(clk), .CD(n18331), .Q(
        poly7_shifted[97]) );
  CFD2QXL \Poly7_reg[102]  ( .D(n10002), .CP(clk), .CD(n18332), .Q(
        poly7_shifted[114]) );
  CFD2QXL \Poly7_reg[159]  ( .D(n9945), .CP(clk), .CD(n18334), .Q(
        poly7_shifted[171]) );
  CFD2QXL \Poly7_reg[164]  ( .D(n9940), .CP(clk), .CD(n18335), .Q(
        poly7_shifted[176]) );
  CFD2QXL \Poly7_reg[224]  ( .D(n9880), .CP(clk), .CD(n18338), .Q(
        poly7_shifted[236]) );
  CFD2QXL \Poly15_reg[1]  ( .D(n9636), .CP(clk), .CD(n18345), .Q(
        poly15_shifted[16]) );
  CFD2QXL \Poly15_reg[3]  ( .D(n9634), .CP(clk), .CD(n18346), .Q(
        poly15_shifted[18]) );
  CFD2QXL \Poly15_reg[2]  ( .D(n9635), .CP(clk), .CD(n18256), .Q(
        poly15_shifted[17]) );
  CFD2QXL \Poly0_reg[90]  ( .D(n9487), .CP(clk), .CD(n18347), .Q(
        poly0_shifted[108]) );
  CFD2QXL \Poly0_reg[80]  ( .D(n9497), .CP(clk), .CD(n18350), .Q(
        poly0_shifted[98]) );
  CFD2QXL \Poly0_reg[79]  ( .D(n9498), .CP(clk), .CD(n18351), .Q(
        poly0_shifted[97]) );
  CFD2QXL \Poly0_reg[84]  ( .D(n9493), .CP(clk), .CD(n18352), .Q(
        poly0_shifted[102]) );
  CFD2QXL \Poly0_reg[81]  ( .D(n9496), .CP(clk), .CD(n18352), .Q(
        poly0_shifted[99]) );
  CFD2QXL \Poly0_reg[86]  ( .D(n9491), .CP(clk), .CD(n18353), .Q(
        poly0_shifted[104]) );
  CFD2QXL \Poly0_reg[83]  ( .D(n9494), .CP(clk), .CD(n18353), .Q(
        poly0_shifted[101]) );
  CFD2QXL \Poly0_reg[88]  ( .D(n9489), .CP(clk), .CD(n18353), .Q(
        poly0_shifted[106]) );
  CFD2QXL \Poly0_reg[78]  ( .D(n9499), .CP(clk), .CD(n18357), .Q(
        poly0_shifted[96]) );
  CFD2QXL \Poly1_reg[305]  ( .D(n9052), .CP(clk), .CD(n18362), .Q(
        poly1_shifted[316]) );
  CFD2QXL \Poly1_reg[145]  ( .D(n9212), .CP(clk), .CD(n18363), .Q(
        poly1_shifted[156]) );
  CFD2QXL \Poly1_reg[189]  ( .D(n9168), .CP(clk), .CD(n18364), .Q(
        poly1_shifted[200]) );
  CFD2QXL \Poly1_reg[177]  ( .D(n9180), .CP(clk), .CD(n18365), .Q(
        poly1_shifted[188]) );
  CFD2QXL \Poly1_reg[247]  ( .D(n9110), .CP(clk), .CD(n18254), .Q(
        poly1_shifted[258]) );
  CFD2QXL \Poly1_reg[313]  ( .D(n9044), .CP(clk), .CD(n18366), .Q(
        poly1_shifted[324]) );
  CFD2QXL \Poly1_reg[131]  ( .D(n9226), .CP(clk), .CD(n18367), .Q(
        poly1_shifted[142]) );
  CFD2QXL \Poly1_reg[174]  ( .D(n9183), .CP(clk), .CD(n18369), .Q(
        poly1_shifted[185]) );
  CFD2QXL \Poly1_reg[96]  ( .D(n9261), .CP(clk), .CD(n18370), .Q(
        poly1_shifted[107]) );
  CFD2QXL \Poly1_reg[255]  ( .D(n9102), .CP(clk), .CD(n18371), .Q(
        poly1_shifted[266]) );
  CFD2QXL \Poly1_reg[265]  ( .D(n9092), .CP(clk), .CD(n18374), .Q(
        poly1_shifted[276]) );
  CFD2QXL \Poly1_reg[127]  ( .D(n9230), .CP(clk), .CD(n18375), .Q(
        poly1_shifted[138]) );
  CFD2QXL \Poly1_reg[81]  ( .D(n9276), .CP(clk), .CD(n18376), .Q(
        poly1_shifted[92]) );
  CFD2QXL \Poly2_reg[7]  ( .D(n9003), .CP(clk), .CD(n18377), .Q(
        poly2_shifted[19]) );
  CFD2QXL \Poly2_reg[3]  ( .D(n9007), .CP(clk), .CD(n18379), .Q(
        poly2_shifted[15]) );
  CFD2QXL \Poly3_reg[20]  ( .D(n8920), .CP(clk), .CD(n18381), .Q(
        poly3_shifted[34]) );
  CFD2QXL \Poly3_reg[23]  ( .D(n8917), .CP(clk), .CD(n18381), .Q(
        poly3_shifted[37]) );
  CFD2QXL \Poly3_reg[12]  ( .D(n8928), .CP(clk), .CD(n18381), .Q(
        poly3_shifted[26]) );
  CFD2QXL \Poly3_reg[15]  ( .D(n8925), .CP(clk), .CD(n18382), .Q(
        poly3_shifted[29]) );
  CFD2QXL \Poly3_reg[27]  ( .D(n8913), .CP(clk), .CD(n18383), .Q(
        poly3_shifted[41]) );
  CFD2QXL \Poly9_reg[47]  ( .D(n11258), .CP(clk), .CD(n18257), .Q(
        poly9_shifted[58]) );
  CFD2QXL \Poly9_reg[75]  ( .D(n11230), .CP(clk), .CD(n18257), .Q(
        poly9_shifted[86]) );
  CFD2QXL \Poly13_reg[60]  ( .D(n11000), .CP(clk), .CD(n18266), .Q(
        poly13_shifted[74]) );
  CFD2QXL \Poly13_reg[211]  ( .D(n10849), .CP(clk), .CD(n18272), .Q(
        poly13_shifted[225]) );
  CFD2QXL \Poly13_reg[497]  ( .D(n10563), .CP(clk), .CD(n18277), .Q(
        poly13_shifted[511]) );
  CFD2QXL \Poly13_reg[250]  ( .D(n10810), .CP(clk), .CD(n18278), .Q(
        poly13_shifted[264]) );
  CFD2QXL \Poly13_reg[423]  ( .D(n10637), .CP(clk), .CD(n18284), .Q(
        poly13_shifted[437]) );
  CFD2QXL \Poly13_reg[437]  ( .D(n10623), .CP(clk), .CD(n18284), .Q(
        poly13_shifted[451]) );
  CFD2QXL \Poly13_reg[451]  ( .D(n10609), .CP(clk), .CD(n18284), .Q(
        poly13_shifted[465]) );
  CFD2QXL \Poly13_reg[329]  ( .D(n10731), .CP(clk), .CD(n18288), .Q(
        poly13_shifted[343]) );
  CFD2QXL \Poly13_reg[343]  ( .D(n10717), .CP(clk), .CD(n18288), .Q(
        poly13_shifted[357]) );
  CFD2QXL \Poly13_reg[357]  ( .D(n10703), .CP(clk), .CD(n18288), .Q(
        poly13_shifted[371]) );
  CFD2QXL \Poly13_reg[371]  ( .D(n10689), .CP(clk), .CD(n18288), .Q(
        poly13_shifted[385]) );
  CFD2QXL \Poly13_reg[303]  ( .D(n10757), .CP(clk), .CD(n18289), .Q(
        poly13_shifted[317]) );
  CFD2QXL \Poly13_reg[317]  ( .D(n10743), .CP(clk), .CD(n18289), .Q(
        poly13_shifted[331]) );
  CFD2QXL \Poly13_reg[331]  ( .D(n10729), .CP(clk), .CD(n18289), .Q(
        poly13_shifted[345]) );
  CFD2QXL \Poly13_reg[345]  ( .D(n10715), .CP(clk), .CD(n18289), .Q(
        poly13_shifted[359]) );
  CFD2QXL \Poly14_reg[240]  ( .D(n10165), .CP(clk), .CD(n18254), .Q(
        poly14_shifted[256]) );
  CFD2QXL \Poly14_reg[67]  ( .D(n10338), .CP(clk), .CD(n18300), .Q(
        poly14_shifted[83]) );
  CFD2QXL \Poly14_reg[109]  ( .D(n10296), .CP(clk), .CD(n18301), .Q(
        poly14_shifted[125]) );
  CFD2QXL \Poly14_reg[10]  ( .D(n10395), .CP(clk), .CD(n18310), .Q(
        poly14_shifted[26]) );
  CFD2QXL \Poly14_reg[106]  ( .D(n10299), .CP(clk), .CD(n18311), .Q(
        poly14_shifted[122]) );
  CFD2QXL \Poly7_reg[231]  ( .D(n9873), .CP(clk), .CD(n18341), .Q(
        poly7_shifted[243]) );
  CFD2QXL \Poly0_reg[2]  ( .D(n9575), .CP(clk), .CD(n18348), .Q(
        poly0_shifted[20]) );
  CFD2QXL \Poly1_reg[121]  ( .D(n9236), .CP(clk), .CD(n18359), .Q(
        poly1_shifted[132]) );
  CFD2QXL \Poly1_reg[308]  ( .D(n9049), .CP(clk), .CD(n18360), .Q(
        poly1_shifted[319]) );
  CFD2QXL \Poly1_reg[252]  ( .D(n9105), .CP(clk), .CD(n18360), .Q(
        poly1_shifted[263]) );
  CFD2QXL \Poly1_reg[285]  ( .D(n9072), .CP(clk), .CD(n18360), .Q(
        poly1_shifted[296]) );
  CFD2QXL \Poly1_reg[173]  ( .D(n9184), .CP(clk), .CD(n18370), .Q(
        poly1_shifted[184]) );
  CFD2QXL \Poly1_reg[288]  ( .D(n9069), .CP(clk), .CD(n18371), .Q(
        poly1_shifted[299]) );
  CFD2QXL \Poly11_reg[45]  ( .D(n11144), .CP(clk), .CD(n18257), .Q(Poly11[45])
         );
  CFD2QXL \Poly11_reg[51]  ( .D(n11138), .CP(clk), .CD(n18257), .Q(Poly11[51])
         );
  CFD2QXL \Poly11_reg[52]  ( .D(n11137), .CP(clk), .CD(n18257), .Q(Poly11[52])
         );
  CFD2QXL \Poly11_reg[42]  ( .D(n11147), .CP(clk), .CD(n18262), .Q(Poly11[42])
         );
  CFD2QXL \Poly7_reg[48]  ( .D(n10056), .CP(clk), .CD(n18316), .Q(Poly7[48])
         );
  CFD2QXL \Poly1_reg[53]  ( .D(n9304), .CP(clk), .CD(n18368), .Q(Poly1[53]) );
  CFD2QXL \Poly4_reg[17]  ( .D(n8839), .CP(clk), .CD(n18384), .Q(Poly4[17]) );
  CFD2QXL \Poly5_reg[96]  ( .D(n11430), .CP(clk), .CD(n18257), .Q(Poly5[96])
         );
  CFD2QXL \Poly8_reg[78]  ( .D(n11323), .CP(clk), .CD(n18257), .Q(Poly8[78])
         );
  CFD2QXL \Poly9_reg[88]  ( .D(n11217), .CP(clk), .CD(n18257), .Q(Poly9[88])
         );
  CFD2QXL \Poly9_reg[87]  ( .D(n11218), .CP(clk), .CD(n18257), .Q(Poly9[87])
         );
  CFD2QXL \Poly9_reg[84]  ( .D(n11221), .CP(clk), .CD(n18257), .Q(Poly9[84])
         );
  CFD2QXL \Poly9_reg[85]  ( .D(n11220), .CP(clk), .CD(n18257), .Q(Poly9[85])
         );
  CFD2QXL \Poly9_reg[86]  ( .D(n11219), .CP(clk), .CD(n18257), .Q(Poly9[86])
         );
  CFD2QXL \Poly11_reg[56]  ( .D(n11133), .CP(clk), .CD(n18257), .Q(Poly11[56])
         );
  CFD2QXL \Poly13_reg[392]  ( .D(n10668), .CP(clk), .CD(n18266), .Q(
        Poly13[392]) );
  CFD2QXL \Poly13_reg[158]  ( .D(n10902), .CP(clk), .CD(n18267), .Q(
        Poly13[158]) );
  CFD2QXL \Poly13_reg[157]  ( .D(n10903), .CP(clk), .CD(n18268), .Q(
        Poly13[157]) );
  CFD2QXL \Poly13_reg[270]  ( .D(n10790), .CP(clk), .CD(n18269), .Q(
        Poly13[270]) );
  CFD2QXL \Poly13_reg[155]  ( .D(n10905), .CP(clk), .CD(n18271), .Q(
        Poly13[155]) );
  CFD2QXL \Poly13_reg[396]  ( .D(n10664), .CP(clk), .CD(n18272), .Q(
        Poly13[396]) );
  CFD2QXL \Poly13_reg[281]  ( .D(n10779), .CP(clk), .CD(n18273), .Q(
        Poly13[281]) );
  CFD2QXL \Poly13_reg[395]  ( .D(n10665), .CP(clk), .CD(n18273), .Q(
        Poly13[395]) );
  CFD2QXL \Poly13_reg[393]  ( .D(n10667), .CP(clk), .CD(n18255), .Q(
        Poly13[393]) );
  CFD2QXL \Poly13_reg[164]  ( .D(n10896), .CP(clk), .CD(n18279), .Q(
        Poly13[164]) );
  CFD2QXL \Poly13_reg[277]  ( .D(n10783), .CP(clk), .CD(n18280), .Q(
        Poly13[277]) );
  CFD2QXL \Poly13_reg[163]  ( .D(n10897), .CP(clk), .CD(n18282), .Q(
        Poly13[163]) );
  CFD2QXL \Poly13_reg[162]  ( .D(n10898), .CP(clk), .CD(n18255), .Q(
        Poly13[162]) );
  CFD2QXL \Poly13_reg[161]  ( .D(n10899), .CP(clk), .CD(n18285), .Q(
        Poly13[161]) );
  CFD2QXL \Poly13_reg[273]  ( .D(n10787), .CP(clk), .CD(n18288), .Q(
        Poly13[273]) );
  CFD2QXL \Poly13_reg[387]  ( .D(n10673), .CP(clk), .CD(n18289), .Q(
        Poly13[387]) );
  CFD2QXL \Poly13_reg[398]  ( .D(n10662), .CP(clk), .CD(n18291), .Q(
        Poly13[398]) );
  CFD2QXL \Poly12_reg[96]  ( .D(n10436), .CP(clk), .CD(n18292), .Q(Poly12[96])
         );
  CFD2QXL \Poly12_reg[19]  ( .D(n10513), .CP(clk), .CD(n18293), .Q(Poly12[19])
         );
  CFD2QXL \Poly12_reg[83]  ( .D(n10449), .CP(clk), .CD(n18294), .Q(Poly12[83])
         );
  CFD2QXL \Poly12_reg[51]  ( .D(n10481), .CP(clk), .CD(n18294), .Q(Poly12[51])
         );
  CFD2QXL \Poly12_reg[87]  ( .D(n10445), .CP(clk), .CD(n18295), .Q(Poly12[87])
         );
  CFD2QXL \Poly12_reg[18]  ( .D(n10514), .CP(clk), .CD(n18298), .Q(Poly12[18])
         );
  CFD2QXL \Poly12_reg[88]  ( .D(n10444), .CP(clk), .CD(n18299), .Q(Poly12[88])
         );
  CFD2QXL \Poly12_reg[86]  ( .D(n10446), .CP(clk), .CD(n18299), .Q(Poly12[86])
         );
  CFD2QXL \Poly14_reg[176]  ( .D(n10229), .CP(clk), .CD(n18254), .Q(
        Poly14[176]) );
  CFD2QXL \Poly14_reg[179]  ( .D(n10226), .CP(clk), .CD(n18300), .Q(
        Poly14[179]) );
  CFD2QXL \Poly14_reg[172]  ( .D(n10233), .CP(clk), .CD(n18308), .Q(
        Poly14[172]) );
  CFD2QXL \Poly14_reg[170]  ( .D(n10235), .CP(clk), .CD(n18311), .Q(
        Poly14[170]) );
  CFD2QXL \Poly14_reg[213]  ( .D(n10192), .CP(clk), .CD(n18312), .Q(
        Poly14[213]) );
  CFD2QXL \Poly14_reg[211]  ( .D(n10194), .CP(clk), .CD(n18316), .Q(
        Poly14[211]) );
  CFD2QXL \Poly7_reg[24]  ( .D(n10080), .CP(clk), .CD(n18316), .Q(Poly7[24])
         );
  CFD2QXL \Poly7_reg[240]  ( .D(n9864), .CP(clk), .CD(n18317), .Q(Poly7[240])
         );
  CFD2QXL \Poly7_reg[21]  ( .D(n10083), .CP(clk), .CD(n18318), .Q(Poly7[21])
         );
  CFD2QXL \Poly7_reg[23]  ( .D(n10081), .CP(clk), .CD(n18319), .Q(Poly7[23])
         );
  CFD2QXL \Poly7_reg[27]  ( .D(n10077), .CP(clk), .CD(n18321), .Q(Poly7[27])
         );
  CFD2QXL \Poly7_reg[29]  ( .D(n10075), .CP(clk), .CD(n18322), .Q(Poly7[29])
         );
  CFD2QXL \Poly7_reg[26]  ( .D(n10078), .CP(clk), .CD(n18325), .Q(Poly7[26])
         );
  CFD2QXL \Poly7_reg[50]  ( .D(n10054), .CP(clk), .CD(n18325), .Q(Poly7[50])
         );
  CFD2QXL \Poly7_reg[57]  ( .D(n10047), .CP(clk), .CD(n18325), .Q(Poly7[57])
         );
  CFD2QXL \Poly7_reg[182]  ( .D(n9922), .CP(clk), .CD(n18326), .Q(Poly7[182])
         );
  CFD2QXL \Poly7_reg[28]  ( .D(n10076), .CP(clk), .CD(n18327), .Q(Poly7[28])
         );
  CFD2QXL \Poly7_reg[59]  ( .D(n10045), .CP(clk), .CD(n18328), .Q(Poly7[59])
         );
  CFD2QXL \Poly7_reg[179]  ( .D(n9925), .CP(clk), .CD(n18328), .Q(Poly7[179])
         );
  CFD2QXL \Poly7_reg[242]  ( .D(n9862), .CP(clk), .CD(n18329), .Q(Poly7[242])
         );
  CFD2QXL \Poly7_reg[30]  ( .D(n10074), .CP(clk), .CD(n18330), .Q(Poly7[30])
         );
  CFD2QXL \Poly7_reg[54]  ( .D(n10050), .CP(clk), .CD(n18331), .Q(Poly7[54])
         );
  CFD2QXL \Poly7_reg[181]  ( .D(n9923), .CP(clk), .CD(n18331), .Q(Poly7[181])
         );
  CFD2QXL \Poly7_reg[244]  ( .D(n9860), .CP(clk), .CD(n18332), .Q(Poly7[244])
         );
  CFD2QXL \Poly7_reg[237]  ( .D(n9867), .CP(clk), .CD(n18333), .Q(Poly7[237])
         );
  CFD2QXL \Poly7_reg[20]  ( .D(n10084), .CP(clk), .CD(n18334), .Q(Poly7[20])
         );
  CFD2QXL \Poly7_reg[56]  ( .D(n10048), .CP(clk), .CD(n18334), .Q(Poly7[56])
         );
  CFD2QXL \Poly7_reg[51]  ( .D(n10053), .CP(clk), .CD(n18334), .Q(Poly7[51])
         );
  CFD2QXL \Poly7_reg[22]  ( .D(n10082), .CP(clk), .CD(n18337), .Q(Poly7[22])
         );
  CFD2QXL \Poly7_reg[53]  ( .D(n10051), .CP(clk), .CD(n18337), .Q(Poly7[53])
         );
  CFD2QXL \Poly7_reg[236]  ( .D(n9868), .CP(clk), .CD(n18338), .Q(Poly7[236])
         );
  CFD2QXL \Poly7_reg[235]  ( .D(n9869), .CP(clk), .CD(n18341), .Q(Poly7[235])
         );
  CFD2QXL \Poly7_reg[238]  ( .D(n9866), .CP(clk), .CD(n18341), .Q(Poly7[238])
         );
  CFD2QXL \Poly0_reg[20]  ( .D(n9557), .CP(clk), .CD(n18348), .Q(Poly0[20]) );
  CFD2QXL \Poly0_reg[10]  ( .D(n9567), .CP(clk), .CD(n18349), .Q(Poly0[10]) );
  CFD2QXL \Poly0_reg[151]  ( .D(n9426), .CP(clk), .CD(n18349), .Q(Poly0[151])
         );
  CFD2QXL \Poly0_reg[150]  ( .D(n9427), .CP(clk), .CD(n18358), .Q(Poly0[150])
         );
  CFD2QXL \Poly1_reg[198]  ( .D(n9159), .CP(clk), .CD(n18359), .Q(Poly1[198])
         );
  CFD2QXL \Poly1_reg[231]  ( .D(n9126), .CP(clk), .CD(n18359), .Q(Poly1[231])
         );
  CFD2QXL \Poly1_reg[157]  ( .D(n9200), .CP(clk), .CD(n18362), .Q(Poly1[157])
         );
  CFD2QXL \Poly1_reg[57]  ( .D(n9300), .CP(clk), .CD(n18363), .Q(Poly1[57]) );
  CFD2QXL \Poly1_reg[156]  ( .D(n9201), .CP(clk), .CD(n18363), .Q(Poly1[156])
         );
  CFD2QXL \Poly1_reg[200]  ( .D(n9157), .CP(clk), .CD(n18364), .Q(Poly1[200])
         );
  CFD2QXL \Poly1_reg[233]  ( .D(n9124), .CP(clk), .CD(n18364), .Q(Poly1[233])
         );
  CFD2QXL \Poly1_reg[155]  ( .D(n9202), .CP(clk), .CD(n18365), .Q(Poly1[155])
         );
  CFD2QXL \Poly1_reg[199]  ( .D(n9158), .CP(clk), .CD(n18254), .Q(Poly1[199])
         );
  CFD2QXL \Poly1_reg[232]  ( .D(n9125), .CP(clk), .CD(n18254), .Q(Poly1[232])
         );
  CFD2QXL \Poly1_reg[54]  ( .D(n9303), .CP(clk), .CD(n18366), .Q(Poly1[54]) );
  CFD2QXL \Poly1_reg[153]  ( .D(n9204), .CP(clk), .CD(n18367), .Q(Poly1[153])
         );
  CFD2QXL \Poly1_reg[230]  ( .D(n9127), .CP(clk), .CD(n18367), .Q(Poly1[230])
         );
  CFD2QXL \Poly1_reg[152]  ( .D(n9205), .CP(clk), .CD(n18369), .Q(Poly1[152])
         );
  CFD2QXL \Poly1_reg[207]  ( .D(n9150), .CP(clk), .CD(n18369), .Q(Poly1[207])
         );
  CFD2QXL \Poly1_reg[229]  ( .D(n9128), .CP(clk), .CD(n18369), .Q(Poly1[229])
         );
  CFD2QXL \Poly1_reg[63]  ( .D(n9294), .CP(clk), .CD(n18370), .Q(Poly1[63]) );
  CFD2QXL \Poly1_reg[151]  ( .D(n9206), .CP(clk), .CD(n18370), .Q(Poly1[151])
         );
  CFD2QXL \Poly1_reg[206]  ( .D(n9151), .CP(clk), .CD(n18371), .Q(Poly1[206])
         );
  CFD2QXL \Poly1_reg[161]  ( .D(n9196), .CP(clk), .CD(n18372), .Q(Poly1[161])
         );
  CFD2QXL \Poly1_reg[205]  ( .D(n9152), .CP(clk), .CD(n18372), .Q(Poly1[205])
         );
  CFD2QXL \Poly1_reg[60]  ( .D(n9297), .CP(clk), .CD(n18373), .Q(Poly1[60]) );
  CFD2QXL \Poly1_reg[159]  ( .D(n9198), .CP(clk), .CD(n18373), .Q(Poly1[159])
         );
  CFD2QXL \Poly1_reg[203]  ( .D(n9154), .CP(clk), .CD(n18373), .Q(Poly1[203])
         );
  CFD2QXL \Poly1_reg[225]  ( .D(n9132), .CP(clk), .CD(n18374), .Q(Poly1[225])
         );
  CFD2QXL \Poly1_reg[227]  ( .D(n9130), .CP(clk), .CD(n18374), .Q(Poly1[227])
         );
  CFD2QXL \Poly1_reg[204]  ( .D(n9153), .CP(clk), .CD(n18375), .Q(Poly1[204])
         );
  CFD2QXL \Poly1_reg[59]  ( .D(n9298), .CP(clk), .CD(n18375), .Q(Poly1[59]) );
  CFD2QXL \Poly1_reg[158]  ( .D(n9199), .CP(clk), .CD(n18376), .Q(Poly1[158])
         );
  CFD2QXL \Poly1_reg[202]  ( .D(n9155), .CP(clk), .CD(n18376), .Q(Poly1[202])
         );
  CFD2QXL \Poly1_reg[235]  ( .D(n9122), .CP(clk), .CD(n18376), .Q(Poly1[235])
         );
  CFD2QXL \Poly1_reg[234]  ( .D(n9123), .CP(clk), .CD(n18377), .Q(Poly1[234])
         );
  CFD2QXL \Poly1_reg[226]  ( .D(n9131), .CP(clk), .CD(n18377), .Q(Poly1[226])
         );
  CFD2QXL \Poly3_reg[34]  ( .D(n8906), .CP(clk), .CD(n18381), .Q(Poly3[34]) );
  CFD2QXL \Poly3_reg[35]  ( .D(n8905), .CP(clk), .CD(n18382), .Q(Poly3[35]) );
  CFD2QXL \Poly3_reg[52]  ( .D(n8888), .CP(clk), .CD(n18383), .Q(Poly3[52]) );
  CFD2QXL \Poly3_reg[33]  ( .D(n8907), .CP(clk), .CD(n18384), .Q(Poly3[33]) );
  CFD2QXL \Poly4_reg[24]  ( .D(n8832), .CP(clk), .CD(n18385), .Q(Poly4[24]) );
  CFD2QXL \Poly4_reg[27]  ( .D(n8829), .CP(clk), .CD(n18386), .Q(Poly4[27]) );
  CFD2QXL \Poly4_reg[3]  ( .D(n8853), .CP(clk), .CD(n18256), .Q(
        poly4_shifted[20]) );
  CFD2QXL \Poly0_reg[103]  ( .D(n9474), .CP(clk), .CD(n18354), .Q(Poly0[103])
         );
  CFD2QXL \Poly0_reg[105]  ( .D(n9472), .CP(clk), .CD(n18355), .Q(Poly0[105])
         );
  CFD2QXL \Poly0_reg[114]  ( .D(n9463), .CP(clk), .CD(n18358), .Q(Poly0[114])
         );
  CFD2QXL \Poly5_reg[28]  ( .D(n11498), .CP(clk), .CD(n18257), .Q(
        poly5_shifted[42]) );
  CFD2QXL \Poly5_reg[27]  ( .D(n11499), .CP(clk), .CD(n18259), .Q(
        poly5_shifted[41]) );
  CFD2QXL \Poly5_reg[41]  ( .D(n11485), .CP(clk), .CD(n18259), .Q(
        poly5_shifted[55]) );
  CFD2QXL \Poly5_reg[59]  ( .D(n11467), .CP(clk), .CD(n18257), .Q(
        poly5_shifted[73]) );
  CFD2QXL \Poly0_reg[91]  ( .D(n9486), .CP(clk), .CD(n18357), .Q(
        poly0_shifted[109]) );
  CFD2QXL \Poly0_reg[113]  ( .D(n9464), .CP(clk), .CD(n18351), .Q(Poly0[113])
         );
  CFD2QXL \Poly0_reg[112]  ( .D(n9465), .CP(clk), .CD(n18356), .Q(Poly0[112])
         );
  CFD2QXL \dataselector_reg[38]  ( .D(n8757), .CP(clk), .CD(n18387), .Q(
        dataselector[38]) );
  CFD2QXL \Poly0_reg[6]  ( .D(n9571), .CP(clk), .CD(n18348), .Q(Poly0[6]) );
  CFD2QXL \scrambler_reg[10]  ( .D(n8710), .CP(clk), .CD(n18257), .Q(
        scrambler[10]) );
  CFD2QXL \Poly15_reg[4]  ( .D(n9633), .CP(clk), .CD(n18345), .Q(
        poly15_shifted[19]) );
  CFD2QXL \Poly5_reg[1]  ( .D(n11525), .CP(clk), .CD(n18257), .Q(Poly5[1]) );
  CFD2QXL \Poly5_reg[2]  ( .D(n11524), .CP(clk), .CD(n18258), .Q(Poly5[2]) );
  CFD2QXL \Poly6_reg[32]  ( .D(n9661), .CP(clk), .CD(n18343), .Q(Poly6[32]) );
  CFD2QXL \dataselector_reg[54]  ( .D(n8741), .CP(clk), .CD(n18257), .Q(
        dataselector[54]) );
  CFD2QXL \Poly6_reg[44]  ( .D(n9649), .CP(clk), .CD(n18344), .Q(Poly6[44]) );
  CFD2QXL \Poly10_reg[7]  ( .D(n11096), .CP(clk), .CD(n18257), .Q(
        poly10_shifted[19]) );
  CFD2QXL \Poly10_reg[3]  ( .D(n11100), .CP(clk), .CD(n18400), .Q(Poly10[3])
         );
  CFD2QXL \dataselector_reg[52]  ( .D(n8743), .CP(clk), .CD(n18402), .Q(
        dataselector[52]) );
  CFD2QXL \Poly10_reg[12]  ( .D(n11091), .CP(clk), .CD(n18262), .Q(Poly10[12])
         );
  CFD2QXL \Poly0_reg[9]  ( .D(n9568), .CP(clk), .CD(n18352), .Q(Poly0[9]) );
  CFD2QXL \Poly3_reg[60]  ( .D(n8880), .CP(clk), .CD(n18390), .Q(
        poly3_shifted[74]) );
  CFD2QXL \Poly13_reg[11]  ( .D(n11049), .CP(clk), .CD(n18277), .Q(
        poly13_shifted[25]) );
  CFD2QXL \dataselector_reg[12]  ( .D(n8783), .CP(clk), .CD(n18388), .Q(
        dataselector[12]) );
  CFD2QXL \Poly12_reg[94]  ( .D(n10438), .CP(clk), .CD(n18297), .Q(Poly12[94])
         );
  CFD2QXL \Poly15_reg[46]  ( .D(n9591), .CP(clk), .CD(n18345), .Q(Poly15[46])
         );
  CFD2QXL \Poly0_reg[119]  ( .D(n9458), .CP(clk), .CD(n18394), .Q(Poly0[119])
         );
  CFD2QXL \Poly0_reg[52]  ( .D(n9525), .CP(clk), .CD(n18395), .Q(
        poly0_shifted[70]) );
  CFD2QXL \Poly10_reg[2]  ( .D(n11101), .CP(clk), .CD(n18263), .Q(Poly10[2])
         );
  CFD2QXL \Poly12_reg[38]  ( .D(n10494), .CP(clk), .CD(n18298), .Q(
        poly12_shifted[54]) );
  CFD2QXL \dataselector_reg[3]  ( .D(n8792), .CP(clk), .CD(n18388), .Q(
        dataselector[3]) );
  CFD2QXL \Poly10_reg[5]  ( .D(n11098), .CP(clk), .CD(n18400), .Q(
        poly10_shifted[17]) );
  CFD2QXL \Poly1_reg[166]  ( .D(n9191), .CP(clk), .CD(n18365), .Q(
        poly1_shifted[177]) );
  CFD2QXL \Poly3_reg[49]  ( .D(n8891), .CP(clk), .CD(n18382), .Q(Poly3[49]) );
  CFD2QXL \Poly1_reg[70]  ( .D(n9287), .CP(clk), .CD(n18376), .Q(
        poly1_shifted[81]) );
  CFD2QXL \Poly11_reg[63]  ( .D(n11126), .CP(clk), .CD(n18257), .Q(Poly11[63])
         );
  CFD2QXL \Poly2_reg[46]  ( .D(n8964), .CP(clk), .CD(n18379), .Q(Poly2[46]) );
  CFD2QXL \Poly4_reg[34]  ( .D(n8822), .CP(clk), .CD(n18384), .Q(Poly4[34]) );
  CFD2QXL \Poly5_reg[95]  ( .D(n11431), .CP(clk), .CD(n18257), .Q(Poly5[95])
         );
  CFD2QXL \Poly12_reg[64]  ( .D(n10468), .CP(clk), .CD(n18292), .Q(Poly12[64])
         );
  CFD2QXL \Poly2_reg[43]  ( .D(n8967), .CP(clk), .CD(n18257), .Q(
        poly2_shifted[55]) );
  CFD2QXL \Poly5_reg[8]  ( .D(n11518), .CP(clk), .CD(n18259), .Q(
        poly5_shifted[22]) );
  CFD2QXL \Poly5_reg[5]  ( .D(n11521), .CP(clk), .CD(n18257), .Q(
        poly5_shifted[19]) );
  CFD2QXL \Poly5_reg[12]  ( .D(n11514), .CP(clk), .CD(n18257), .Q(
        poly5_shifted[26]) );
  CFD2QXL \Poly8_reg[25]  ( .D(n11376), .CP(clk), .CD(n18261), .Q(
        poly8_shifted[39]) );
  CFD2QXL \Poly8_reg[23]  ( .D(n11378), .CP(clk), .CD(n18257), .Q(
        poly8_shifted[37]) );
  CFD2QXL \Poly10_reg[27]  ( .D(n11076), .CP(clk), .CD(n18400), .Q(
        poly10_shifted[39]) );
  CFD2QXL \Poly10_reg[8]  ( .D(n11095), .CP(clk), .CD(n18400), .Q(
        poly10_shifted[20]) );
  CFD2QXL \Poly14_reg[226]  ( .D(n10179), .CP(clk), .CD(n18304), .Q(
        poly14_shifted[242]) );
  CFD2QXL \Poly1_reg[244]  ( .D(n9113), .CP(clk), .CD(n18371), .Q(
        poly1_shifted[255]) );
  CFD2QXL \Poly4_reg[12]  ( .D(n8844), .CP(clk), .CD(n18385), .Q(
        poly4_shifted[29]) );
  CFD2QXL \Poly10_reg[28]  ( .D(n11075), .CP(clk), .CD(n18264), .Q(
        poly10_shifted[40]) );
  CFD2QXL \Poly7_reg[40]  ( .D(n10064), .CP(clk), .CD(n18327), .Q(
        poly7_shifted[52]) );
  CFD2QXL \Poly15_reg[35]  ( .D(n9602), .CP(clk), .CD(n18346), .Q(
        poly15_shifted[50]) );
  CFD2QXL \Poly1_reg[163]  ( .D(n9194), .CP(clk), .CD(n18369), .Q(
        poly1_shifted[174]) );
  CFD2QXL \Poly4_reg[8]  ( .D(n8848), .CP(clk), .CD(n18256), .Q(
        poly4_shifted[25]) );
  CFD2QXL \Poly12_reg[110]  ( .D(n10422), .CP(clk), .CD(n18294), .Q(
        poly12_shifted[126]) );
  CFD2QXL \Poly2_reg[36]  ( .D(n8974), .CP(clk), .CD(n18257), .Q(Poly2[36]) );
  CFD2QXL \Poly11_reg[14]  ( .D(n11175), .CP(clk), .CD(n18257), .Q(
        poly11_shifted[29]) );
  CFD2QXL \Poly11_reg[60]  ( .D(n11129), .CP(clk), .CD(n18257), .Q(Poly11[60])
         );
  CFD2QXL \Poly11_reg[57]  ( .D(n11132), .CP(clk), .CD(n18262), .Q(Poly11[57])
         );
  CFD2QXL \Poly8_reg[17]  ( .D(n11384), .CP(clk), .CD(n18257), .Q(
        poly8_shifted[31]) );
  CFD2QXL \Poly10_reg[6]  ( .D(n11097), .CP(clk), .CD(n18400), .Q(
        poly10_shifted[18]) );
  CFD2QXL \Poly0_reg[22]  ( .D(n9555), .CP(clk), .CD(n18348), .Q(Poly0[22]) );
  CFD2QXL \Poly0_reg[178]  ( .D(n9399), .CP(clk), .CD(n18349), .Q(
        poly0_shifted[196]) );
  CFD2QXL \Poly0_reg[50]  ( .D(n9527), .CP(clk), .CD(n18395), .Q(
        poly0_shifted[68]) );
  CFD2QXL \Poly0_reg[181]  ( .D(n9396), .CP(clk), .CD(n18354), .Q(
        poly0_shifted[199]) );
  CFD2QXL \Poly0_reg[184]  ( .D(n9393), .CP(clk), .CD(n18347), .Q(
        poly0_shifted[202]) );
  CFD2QXL \Poly0_reg[190]  ( .D(n9387), .CP(clk), .CD(n18393), .Q(
        poly0_shifted[208]) );
  CFD2QXL \Poly0_reg[176]  ( .D(n9401), .CP(clk), .CD(n18349), .Q(
        poly0_shifted[194]) );
  CFD2QXL \Poly2_reg[29]  ( .D(n8981), .CP(clk), .CD(n18379), .Q(Poly2[29]) );
  CFD2QXL \Poly7_reg[92]  ( .D(n10012), .CP(clk), .CD(n18335), .Q(
        poly7_shifted[104]) );
  CFD2QXL \dataselector_reg[18]  ( .D(n8777), .CP(clk), .CD(n18402), .Q(
        dataselector[18]) );
  CFD2QXL \Poly9_reg[31]  ( .D(n11274), .CP(clk), .CD(n18257), .Q(
        poly9_shifted[42]) );
  CFD2QXL \Poly10_reg[30]  ( .D(n11073), .CP(clk), .CD(n18264), .Q(
        poly10_shifted[42]) );
  CFD2QXL \Poly12_reg[42]  ( .D(n10490), .CP(clk), .CD(n18296), .Q(
        poly12_shifted[58]) );
  CFD2QXL \Poly12_reg[74]  ( .D(n10458), .CP(clk), .CD(n18296), .Q(
        poly12_shifted[90]) );
  CFD2QXL \Poly7_reg[6]  ( .D(n10098), .CP(clk), .CD(n18330), .Q(
        poly7_shifted[18]) );
  CFD2QXL \Poly7_reg[67]  ( .D(n10037), .CP(clk), .CD(n18340), .Q(
        poly7_shifted[79]) );
  CFD2QXL \Poly1_reg[245]  ( .D(n9112), .CP(clk), .CD(n18369), .Q(
        poly1_shifted[256]) );
  CFD2QXL \Poly4_reg[9]  ( .D(n8847), .CP(clk), .CD(n18385), .Q(
        poly4_shifted[26]) );
  CFD2QXL \Poly11_reg[58]  ( .D(n11131), .CP(clk), .CD(n18257), .Q(Poly11[58])
         );
  CFD2QXL \Poly6_reg[23]  ( .D(n9670), .CP(clk), .CD(n18343), .Q(Poly6[23]) );
  CFD2QXL \Poly6_reg[34]  ( .D(n9659), .CP(clk), .CD(n18344), .Q(Poly6[34]) );
  CFD2QXL \Poly9_reg[97]  ( .D(n11208), .CP(clk), .CD(n18257), .Q(
        poly9_shifted[108]) );
  CFD2QXL \Poly12_reg[7]  ( .D(n10525), .CP(clk), .CD(n18293), .Q(
        poly12_shifted[23]) );
  CFD2QXL \Poly12_reg[72]  ( .D(n10460), .CP(clk), .CD(n18299), .Q(
        poly12_shifted[88]) );
  CFD2QXL \Poly14_reg[192]  ( .D(n10213), .CP(clk), .CD(n18254), .Q(
        poly14_shifted[208]) );
  CFD2QXL \Poly4_reg[14]  ( .D(n8842), .CP(clk), .CD(n18385), .Q(
        poly4_shifted[31]) );
  CFD2QXL \Poly12_reg[97]  ( .D(n10435), .CP(clk), .CD(n18298), .Q(
        poly12_shifted[113]) );
  CFD2QXL \Poly14_reg[59]  ( .D(n10346), .CP(clk), .CD(n18304), .Q(
        poly14_shifted[75]) );
  CFD2QXL \Poly0_reg[34]  ( .D(n9543), .CP(clk), .CD(n18353), .Q(
        poly0_shifted[52]) );
  CFD2QXL \Poly0_reg[31]  ( .D(n9546), .CP(clk), .CD(n18354), .Q(
        poly0_shifted[49]) );
  CFD2QXL \Poly0_reg[128]  ( .D(n9449), .CP(clk), .CD(n18355), .Q(
        poly0_shifted[146]) );
  CFD2QXL \Poly3_reg[69]  ( .D(n8871), .CP(clk), .CD(n18383), .Q(
        poly3_shifted[83]) );
  CFD2QXL \Poly3_reg[67]  ( .D(n8873), .CP(clk), .CD(n18384), .Q(
        poly3_shifted[81]) );
  CFD2QXL \Poly3_reg[63]  ( .D(n8877), .CP(clk), .CD(n18382), .Q(
        poly3_shifted[77]) );
  CFD2QXL \Poly14_reg[35]  ( .D(n10370), .CP(clk), .CD(n18254), .Q(
        poly14_shifted[51]) );
  CFD2QXL \Poly7_reg[367]  ( .D(n9737), .CP(clk), .CD(n18327), .Q(
        poly7_shifted[379]) );
  CFD2QXL \Poly9_reg[41]  ( .D(n11264), .CP(clk), .CD(n18257), .Q(
        poly9_shifted[52]) );
  CFD2QXL \Poly9_reg[42]  ( .D(n11263), .CP(clk), .CD(n18257), .Q(
        poly9_shifted[53]) );
  CFD2QXL \Poly7_reg[73]  ( .D(n10031), .CP(clk), .CD(n18331), .Q(
        poly7_shifted[85]) );
  CFD2QXL \dataselector_reg[11]  ( .D(n8784), .CP(clk), .CD(n18402), .Q(
        dataselector[11]) );
  CFD2QXL \Poly5_reg[10]  ( .D(n11516), .CP(clk), .CD(n18260), .Q(
        poly5_shifted[24]) );
  CFD2QXL \Poly1_reg[71]  ( .D(n9286), .CP(clk), .CD(n18373), .Q(
        poly1_shifted[82]) );
  CFD2QXL \dataselector_reg[13]  ( .D(n8782), .CP(clk), .CD(n18388), .Q(
        dataselector[13]) );
  CFD2QXL \Poly5_reg[77]  ( .D(n11449), .CP(clk), .CD(n18257), .Q(Poly5[77])
         );
  CFD2QXL \Poly5_reg[97]  ( .D(n11429), .CP(clk), .CD(n18257), .Q(Poly5[97])
         );
  CFD2QXL \Poly10_reg[4]  ( .D(n11099), .CP(clk), .CD(n18262), .Q(Poly10[4])
         );
  CFD2QXL \Poly10_reg[16]  ( .D(n11087), .CP(clk), .CD(n18264), .Q(Poly10[16])
         );
  CFD2QXL \Poly12_reg[32]  ( .D(n10500), .CP(clk), .CD(n18292), .Q(Poly12[32])
         );
  CFD2QXL \Poly10_reg[10]  ( .D(n11093), .CP(clk), .CD(n18262), .Q(Poly10[10])
         );
  CFD2QXL \Poly14_reg[194]  ( .D(n10211), .CP(clk), .CD(n18316), .Q(
        Poly14[194]) );
  CFD2QXL \Poly14_reg[210]  ( .D(n10195), .CP(clk), .CD(n18316), .Q(
        Poly14[210]) );
  CFD2QXL \Poly6_reg[21]  ( .D(n9672), .CP(clk), .CD(n18343), .Q(Poly6[21]) );
  CFD2QXL \Poly4_reg[38]  ( .D(n8818), .CP(clk), .CD(n18385), .Q(Poly4[38]) );
  CFD2QXL \Poly4_reg[39]  ( .D(n8817), .CP(clk), .CD(n18389), .Q(Poly4[39]) );
  CFD2QXL \Poly10_reg[13]  ( .D(n11090), .CP(clk), .CD(n18400), .Q(Poly10[13])
         );
  CFD2QXL \Poly13_reg[274]  ( .D(n10786), .CP(clk), .CD(n18286), .Q(
        Poly13[274]) );
  CFD2QXL \Poly5_reg[82]  ( .D(n11444), .CP(clk), .CD(n18257), .Q(Poly5[82])
         );
  CFD2QXL \Poly9_reg[3]  ( .D(n11302), .CP(clk), .CD(n18257), .Q(
        poly9_shifted[14]) );
  CFD2QXL \Poly6_reg[17]  ( .D(n9676), .CP(clk), .CD(n18343), .Q(Poly6[17]) );
  CFD2QXL \Poly5_reg[79]  ( .D(n11447), .CP(clk), .CD(n18260), .Q(Poly5[79])
         );
  CFD2QXL \dataselector_reg[49]  ( .D(n8746), .CP(clk), .CD(n18402), .Q(
        dataselector[49]) );
  CFD2QXL \Poly5_reg[91]  ( .D(n11435), .CP(clk), .CD(n18257), .Q(Poly5[91])
         );
  CFD2QXL \Poly11_reg[34]  ( .D(n11155), .CP(clk), .CD(n18257), .Q(Poly11[34])
         );
  CFD2QXL \Poly11_reg[33]  ( .D(n11156), .CP(clk), .CD(n18257), .Q(Poly11[33])
         );
  CFD2QXL \Poly12_reg[93]  ( .D(n10439), .CP(clk), .CD(n18297), .Q(Poly12[93])
         );
  CFD2QXL \Poly9_reg[89]  ( .D(n11216), .CP(clk), .CD(n18257), .Q(Poly9[89])
         );
  CFD2QXL \Poly3_reg[42]  ( .D(n8898), .CP(clk), .CD(n18380), .Q(Poly3[42]) );
  CFD2QXL \Poly10_reg[18]  ( .D(n11085), .CP(clk), .CD(n18263), .Q(Poly10[18])
         );
  CFD2QXL \Poly2_reg[34]  ( .D(n8976), .CP(clk), .CD(n18391), .Q(Poly2[34]) );
  CFD2QXL \Poly8_reg[44]  ( .D(n11357), .CP(clk), .CD(n18257), .Q(
        poly8_shifted[58]) );
  CFD2QXL \Poly3_reg[22]  ( .D(n8918), .CP(clk), .CD(n18384), .Q(
        poly3_shifted[36]) );
  CFD2QXL \Poly5_reg[20]  ( .D(n11506), .CP(clk), .CD(n18257), .Q(
        poly5_shifted[34]) );
  CFD2QXL \Poly5_reg[68]  ( .D(n11458), .CP(clk), .CD(n18257), .Q(
        poly5_shifted[82]) );
  CFD2QXL \Poly5_reg[43]  ( .D(n11483), .CP(clk), .CD(n18257), .Q(
        poly5_shifted[57]) );
  CFD2QXL \Poly9_reg[49]  ( .D(n11256), .CP(clk), .CD(n18257), .Q(
        poly9_shifted[60]) );
  CFD2QXL \Poly12_reg[46]  ( .D(n10486), .CP(clk), .CD(n18398), .Q(
        poly12_shifted[62]) );
  CFD2QXL \Poly6_reg[8]  ( .D(n9685), .CP(clk), .CD(n18396), .Q(
        poly6_shifted[18]) );
  CFD2QXL \Poly0_reg[200]  ( .D(n9377), .CP(clk), .CD(n18347), .Q(
        poly0_shifted[218]) );
  CFD2QXL \Poly0_reg[194]  ( .D(n9383), .CP(clk), .CD(n18349), .Q(
        poly0_shifted[212]) );
  CFD2QXL \Poly5_reg[35]  ( .D(n11491), .CP(clk), .CD(n18257), .Q(
        poly5_shifted[49]) );
  CFD2QXL \Poly11_reg[23]  ( .D(n11166), .CP(clk), .CD(n18257), .Q(Poly11[23])
         );
  CFD2QXL \Poly2_reg[21]  ( .D(n8989), .CP(clk), .CD(n18391), .Q(Poly2[21]) );
  CFD2QXL \Poly10_reg[15]  ( .D(n11088), .CP(clk), .CD(n18263), .Q(Poly10[15])
         );
  CFD2QXL \Poly12_reg[54]  ( .D(n10478), .CP(clk), .CD(n18298), .Q(Poly12[54])
         );
  CFD2QXL \Poly6_reg[40]  ( .D(n9653), .CP(clk), .CD(n18341), .Q(Poly6[40]) );
  CFD2QXL \Poly6_reg[12]  ( .D(n9681), .CP(clk), .CD(n18343), .Q(Poly6[12]) );
  CFD2QXL \Poly3_reg[32]  ( .D(n8908), .CP(clk), .CD(n18390), .Q(Poly3[32]) );
  CFD2QXL \Poly2_reg[31]  ( .D(n8979), .CP(clk), .CD(n18391), .Q(Poly2[31]) );
  CFD2QXL \Poly1_reg[23]  ( .D(n9334), .CP(clk), .CD(n18365), .Q(Poly1[23]) );
  CFD2QXL \Poly11_reg[50]  ( .D(n11139), .CP(clk), .CD(n18257), .Q(Poly11[50])
         );
  CFD2QXL \Poly11_reg[65]  ( .D(n11124), .CP(clk), .CD(n18257), .Q(Poly11[65])
         );
  CFD2QXL \Poly5_reg[92]  ( .D(n11434), .CP(clk), .CD(n18259), .Q(Poly5[92])
         );
  CFD2QXL \Poly8_reg[75]  ( .D(n11326), .CP(clk), .CD(n18257), .Q(Poly8[75])
         );
  CFD2QXL \Poly9_reg[15]  ( .D(n11290), .CP(clk), .CD(n18257), .Q(Poly9[15])
         );
  CFD2QXL \Poly13_reg[282]  ( .D(n10778), .CP(clk), .CD(n18271), .Q(
        Poly13[282]) );
  CFD2QXL \Poly13_reg[276]  ( .D(n10784), .CP(clk), .CD(n18282), .Q(
        Poly13[276]) );
  CFD2QXL \Poly13_reg[275]  ( .D(n10785), .CP(clk), .CD(n18255), .Q(
        Poly13[275]) );
  CFD2QXL \Poly13_reg[388]  ( .D(n10672), .CP(clk), .CD(n18286), .Q(
        Poly13[388]) );
  CFD2QXL \Poly14_reg[167]  ( .D(n10238), .CP(clk), .CD(n18302), .Q(
        Poly14[167]) );
  CFD2QXL \Poly14_reg[166]  ( .D(n10239), .CP(clk), .CD(n18309), .Q(
        Poly14[166]) );
  CFD2QXL \Poly7_reg[234]  ( .D(n9870), .CP(clk), .CD(n18335), .Q(Poly7[234])
         );
  CFD2QXL \Poly7_reg[243]  ( .D(n9861), .CP(clk), .CD(n18341), .Q(Poly7[243])
         );
  CFD2QXL \Poly1_reg[58]  ( .D(n9299), .CP(clk), .CD(n18362), .Q(Poly1[58]) );
  CFD2QXL \Poly1_reg[62]  ( .D(n9295), .CP(clk), .CD(n18372), .Q(Poly1[62]) );
  CFD2QXL \Poly14_reg[218]  ( .D(n10187), .CP(clk), .CD(n18397), .Q(
        poly14_shifted[234]) );
  CFD2QXL \Poly8_reg[24]  ( .D(n11377), .CP(clk), .CD(n18257), .Q(
        poly8_shifted[38]) );
  CFD2QXL \Poly7_reg[218]  ( .D(n9886), .CP(clk), .CD(n18397), .Q(
        poly7_shifted[230]) );
  CFD2QXL \Poly7_reg[90]  ( .D(n10014), .CP(clk), .CD(n18397), .Q(
        poly7_shifted[102]) );
  CFD2QXL \scrambler_reg[15]  ( .D(n8715), .CP(clk), .CD(n18257), .Q(
        scrambler[15]) );
  CFD2QXL \Poly9_reg[33]  ( .D(n11272), .CP(clk), .CD(n18257), .Q(
        poly9_shifted[44]) );
  CFD2QXL \dataselector_reg[30]  ( .D(n8765), .CP(clk), .CD(n18257), .Q(
        dataselector[30]) );
  CFD2QXL \Poly15_reg[21]  ( .D(n9616), .CP(clk), .CD(n18256), .Q(Poly15[21])
         );
  CFD2QXL \Poly5_reg[22]  ( .D(n11504), .CP(clk), .CD(n18259), .Q(
        poly5_shifted[36]) );
  CFD2QXL \Poly5_reg[62]  ( .D(n11464), .CP(clk), .CD(n18257), .Q(
        poly5_shifted[76]) );
  CFD2QXL \Poly5_reg[38]  ( .D(n11488), .CP(clk), .CD(n18260), .Q(
        poly5_shifted[52]) );
  CFD2QXL \Poly8_reg[58]  ( .D(n11343), .CP(clk), .CD(n18257), .Q(
        poly8_shifted[72]) );
  CFD2QXL \Poly11_reg[24]  ( .D(n11165), .CP(clk), .CD(n18257), .Q(Poly11[24])
         );
  CFD2QXL \Poly8_reg[39]  ( .D(n11362), .CP(clk), .CD(n18261), .Q(
        poly8_shifted[53]) );
  CFD2QXL \Poly0_reg[93]  ( .D(n9484), .CP(clk), .CD(n18350), .Q(
        poly0_shifted[111]) );
  CFD2QXL \Poly2_reg[17]  ( .D(n8993), .CP(clk), .CD(n18379), .Q(
        poly2_shifted[29]) );
  CFD2QXL \Poly11_reg[38]  ( .D(n11151), .CP(clk), .CD(n18257), .Q(Poly11[38])
         );
  CFD2QXL \Poly3_reg[54]  ( .D(n8886), .CP(clk), .CD(n18381), .Q(Poly3[54]) );
  CFD2QXL \Poly5_reg[112]  ( .D(n11414), .CP(clk), .CD(n18257), .Q(Poly5[112])
         );
  CFD2QXL \Poly5_reg[113]  ( .D(n11413), .CP(clk), .CD(n18258), .Q(Poly5[113])
         );
  CFD2QXL \Poly5_reg[117]  ( .D(n11409), .CP(clk), .CD(n18257), .Q(Poly5[117])
         );
  CFD2QXL \Poly6_reg[48]  ( .D(n9645), .CP(clk), .CD(n18342), .Q(Poly6[48]) );
  CFD2QXL \Poly9_reg[60]  ( .D(n11245), .CP(clk), .CD(n18257), .Q(
        poly9_shifted[71]) );
  CFD2QXL \dataselector_reg[42]  ( .D(n8753), .CP(clk), .CD(n18402), .Q(
        dataselector[42]) );
  CFD2QXL \scrambler_reg[14]  ( .D(n8714), .CP(clk), .CD(n18257), .Q(
        scrambler[14]) );
  CFD2QXL \scrambler_reg[5]  ( .D(n8705), .CP(clk), .CD(n18257), .Q(
        scrambler[5]) );
  CFD2QXL \Poly9_reg[38]  ( .D(n11267), .CP(clk), .CD(n18257), .Q(
        poly9_shifted[49]) );
  CFD2QXL \Poly1_reg[294]  ( .D(n9063), .CP(clk), .CD(n18392), .Q(
        poly1_shifted[305]) );
  CFD2QXL \Poly5_reg[44]  ( .D(n11482), .CP(clk), .CD(n18258), .Q(
        poly5_shifted[58]) );
  CFD2QXL \Poly8_reg[3]  ( .D(n11398), .CP(clk), .CD(n18257), .Q(Poly8[3]) );
  CFD2QXL \Poly8_reg[74]  ( .D(n11327), .CP(clk), .CD(n18257), .Q(Poly8[74])
         );
  CFD2QXL \Poly9_reg[23]  ( .D(n11282), .CP(clk), .CD(n18257), .Q(Poly9[23])
         );
  CFD2QXL \Poly9_reg[93]  ( .D(n11212), .CP(clk), .CD(n18257), .Q(Poly9[93])
         );
  CFD2QXL \Poly11_reg[68]  ( .D(n11121), .CP(clk), .CD(n18262), .Q(Poly11[68])
         );
  CFD2QXL \Poly13_reg[394]  ( .D(n10666), .CP(clk), .CD(n18275), .Q(
        Poly13[394]) );
  CFD2QXL \Poly12_reg[27]  ( .D(n10505), .CP(clk), .CD(n18293), .Q(Poly12[27])
         );
  CFD2QXL \Poly15_reg[17]  ( .D(n9620), .CP(clk), .CD(n18256), .Q(Poly15[17])
         );
  CFD2QXL \Poly2_reg[50]  ( .D(n8960), .CP(clk), .CD(n18378), .Q(Poly2[50]) );
  CFD2QXL \Poly2_reg[54]  ( .D(n8956), .CP(clk), .CD(n18378), .Q(Poly2[54]) );
  CFD2QXL \Poly1_reg[134]  ( .D(n9223), .CP(clk), .CD(n18392), .Q(
        poly1_shifted[145]) );
  CFD2QXL \Poly9_reg[22]  ( .D(n11283), .CP(clk), .CD(n18257), .Q(Poly9[22])
         );
  CFD2QXL \Poly9_reg[17]  ( .D(n11288), .CP(clk), .CD(n18257), .Q(Poly9[17])
         );
  CFD2QXL \Poly9_reg[91]  ( .D(n11214), .CP(clk), .CD(n18257), .Q(Poly9[91])
         );
  CFD2QXL \Poly9_reg[94]  ( .D(n11211), .CP(clk), .CD(n18257), .Q(Poly9[94])
         );
  CFD2QXL \Poly11_reg[17]  ( .D(n11172), .CP(clk), .CD(n18257), .Q(Poly11[17])
         );
  CFD2QXL \Poly12_reg[29]  ( .D(n10503), .CP(clk), .CD(n18294), .Q(Poly12[29])
         );
  CFD2QXL \Poly12_reg[58]  ( .D(n10474), .CP(clk), .CD(n18296), .Q(Poly12[58])
         );
  CFD2QXL \Poly12_reg[28]  ( .D(n10504), .CP(clk), .CD(n18296), .Q(Poly12[28])
         );
  CFD2QXL \Poly7_reg[187]  ( .D(n9917), .CP(clk), .CD(n18340), .Q(Poly7[187])
         );
  CFD2QXL \Poly15_reg[12]  ( .D(n9625), .CP(clk), .CD(n18345), .Q(Poly15[12])
         );
  CFD2QXL \Poly3_reg[41]  ( .D(n8899), .CP(clk), .CD(n18383), .Q(Poly3[41]) );
  CFD2QXL \Poly4_reg[32]  ( .D(n8824), .CP(clk), .CD(n18256), .Q(Poly4[32]) );
  CFD2QXL \Poly3_reg[61]  ( .D(n8879), .CP(clk), .CD(n18257), .Q(
        poly3_shifted[75]) );
  CFD2QXL \Poly11_reg[46]  ( .D(n11143), .CP(clk), .CD(n18257), .Q(Poly11[46])
         );
  CFD2QXL \Poly14_reg[205]  ( .D(n10200), .CP(clk), .CD(n18315), .Q(
        Poly14[205]) );
  CFD2QXL \Poly6_reg[19]  ( .D(n9674), .CP(clk), .CD(n18342), .Q(Poly6[19]) );
  CFD2QXL \Poly15_reg[24]  ( .D(n9613), .CP(clk), .CD(n18256), .Q(Poly15[24])
         );
  CFD2QXL \Poly2_reg[24]  ( .D(n8986), .CP(clk), .CD(n18377), .Q(Poly2[24]) );
  CFD2QXL \Poly2_reg[26]  ( .D(n8984), .CP(clk), .CD(n18377), .Q(Poly2[26]) );
  CFD2QXL \Poly4_reg[20]  ( .D(n8836), .CP(clk), .CD(n18256), .Q(Poly4[20]) );
  CFD2QXL \Poly4_reg[22]  ( .D(n8834), .CP(clk), .CD(n18386), .Q(Poly4[22]) );
  CFD2QXL \Poly4_reg[30]  ( .D(n8826), .CP(clk), .CD(n18256), .Q(Poly4[30]) );
  CFD2QXL \Poly4_reg[23]  ( .D(n8833), .CP(clk), .CD(n18256), .Q(Poly4[23]) );
  CFD2QXL \Poly5_reg[74]  ( .D(n11452), .CP(clk), .CD(n18257), .Q(
        poly5_shifted[88]) );
  CFD2QXL \Poly8_reg[33]  ( .D(n11368), .CP(clk), .CD(n18257), .Q(
        poly8_shifted[47]) );
  CFD2QXL \Poly9_reg[78]  ( .D(n11227), .CP(clk), .CD(n18257), .Q(
        poly9_shifted[89]) );
  CFD2QXL \Poly9_reg[68]  ( .D(n11237), .CP(clk), .CD(n18257), .Q(
        poly9_shifted[79]) );
  CFD2QXL \Poly11_reg[9]  ( .D(n11180), .CP(clk), .CD(n18257), .Q(
        poly11_shifted[24]) );
  CFD2QXL \Poly13_reg[140]  ( .D(n10920), .CP(clk), .CD(n18399), .Q(
        poly13_shifted[154]) );
  CFD2QXL \Poly13_reg[72]  ( .D(n10988), .CP(clk), .CD(n18400), .Q(
        poly13_shifted[86]) );
  CFD2QXL \Poly13_reg[241]  ( .D(n10819), .CP(clk), .CD(n18399), .Q(
        poly13_shifted[255]) );
  CFD2QXL \Poly13_reg[113]  ( .D(n10947), .CP(clk), .CD(n18399), .Q(
        poly13_shifted[127]) );
  CFD2QXL \Poly13_reg[96]  ( .D(n10964), .CP(clk), .CD(n18400), .Q(
        poly13_shifted[110]) );
  CFD2QXL \Poly13_reg[351]  ( .D(n10709), .CP(clk), .CD(n18399), .Q(
        poly13_shifted[365]) );
  CFD2QXL \Poly13_reg[151]  ( .D(n10909), .CP(clk), .CD(n18399), .Q(
        poly13_shifted[165]) );
  CFD2QXL \Poly13_reg[481]  ( .D(n10579), .CP(clk), .CD(n18399), .Q(
        poly13_shifted[495]) );
  CFD2QXL \Poly13_reg[479]  ( .D(n10581), .CP(clk), .CD(n18399), .Q(
        poly13_shifted[493]) );
  CFD2QXL \Poly13_reg[436]  ( .D(n10624), .CP(clk), .CD(n18399), .Q(
        poly13_shifted[450]) );
  CFD2QXL \Poly12_reg[0]  ( .D(n10532), .CP(clk), .CD(n18398), .Q(
        poly12_shifted[16]) );
  CFD2QXL \Poly14_reg[49]  ( .D(n10356), .CP(clk), .CD(n18398), .Q(
        poly14_shifted[65]) );
  CFD2QXL \Poly14_reg[57]  ( .D(n10348), .CP(clk), .CD(n18398), .Q(
        poly14_shifted[73]) );
  CFD2QXL \Poly14_reg[153]  ( .D(n10252), .CP(clk), .CD(n18398), .Q(
        poly14_shifted[169]) );
  CFD2QXL \Poly14_reg[102]  ( .D(n10303), .CP(clk), .CD(n18398), .Q(
        poly14_shifted[118]) );
  CFD2QXL \Poly14_reg[62]  ( .D(n10343), .CP(clk), .CD(n18398), .Q(
        poly14_shifted[78]) );
  CFD2QXL \Poly7_reg[278]  ( .D(n9826), .CP(clk), .CD(n18397), .Q(
        poly7_shifted[290]) );
  CFD2QXL \Poly7_reg[147]  ( .D(n9957), .CP(clk), .CD(n18397), .Q(
        poly7_shifted[159]) );
  CFD2QXL \Poly7_reg[152]  ( .D(n9952), .CP(clk), .CD(n18397), .Q(
        poly7_shifted[164]) );
  CFD2QXL \Poly7_reg[46]  ( .D(n10058), .CP(clk), .CD(n18397), .Q(
        poly7_shifted[58]) );
  CFD2QXL \Poly15_reg[10]  ( .D(n9627), .CP(clk), .CD(n18396), .Q(
        poly15_shifted[25]) );
  CFD2QXL \Poly1_reg[178]  ( .D(n9179), .CP(clk), .CD(n18392), .Q(
        poly1_shifted[189]) );
  CFD2QXL \Poly1_reg[85]  ( .D(n9272), .CP(clk), .CD(n18392), .Q(
        poly1_shifted[96]) );
  CFD2QXL \Poly1_reg[254]  ( .D(n9103), .CP(clk), .CD(n18392), .Q(
        poly1_shifted[265]) );
  CFD2QXL \Poly2_reg[13]  ( .D(n8997), .CP(clk), .CD(n18391), .Q(
        poly2_shifted[25]) );
  CFD2QXL \Poly3_reg[28]  ( .D(n8912), .CP(clk), .CD(n18390), .Q(
        poly3_shifted[42]) );
  CFD2QXL \Poly4_reg[2]  ( .D(n8854), .CP(clk), .CD(n18389), .Q(
        poly4_shifted[19]) );
  CFD2QXL \Poly5_reg[11]  ( .D(n11515), .CP(clk), .CD(n18257), .Q(
        poly5_shifted[25]) );
  CFD2QXL \Poly8_reg[30]  ( .D(n11371), .CP(clk), .CD(n18257), .Q(
        poly8_shifted[44]) );
  CFD2QXL \Poly8_reg[36]  ( .D(n11365), .CP(clk), .CD(n18257), .Q(
        poly8_shifted[50]) );
  CFD2QXL \Poly8_reg[20]  ( .D(n11381), .CP(clk), .CD(n18257), .Q(
        poly8_shifted[34]) );
  CFD2QXL \Poly9_reg[100]  ( .D(n11205), .CP(clk), .CD(n18257), .Q(
        poly9_shifted[111]) );
  CFD2QXL \Poly13_reg[418]  ( .D(n10642), .CP(clk), .CD(n18399), .Q(
        poly13_shifted[432]) );
  CFD2QXL \Poly13_reg[338]  ( .D(n10722), .CP(clk), .CD(n18399), .Q(
        poly13_shifted[352]) );
  CFD2QXL \Poly13_reg[411]  ( .D(n10649), .CP(clk), .CD(n18399), .Q(
        poly13_shifted[425]) );
  CFD2QXL \Poly13_reg[299]  ( .D(n10761), .CP(clk), .CD(n18399), .Q(
        poly13_shifted[313]) );
  CFD2QXL \Poly14_reg[248]  ( .D(n10157), .CP(clk), .CD(n18397), .Q(
        poly14_shifted[264]) );
  CFD2QXL \Poly14_reg[155]  ( .D(n10250), .CP(clk), .CD(n18398), .Q(
        poly14_shifted[171]) );
  CFD2QXL \Poly14_reg[117]  ( .D(n10288), .CP(clk), .CD(n18398), .Q(
        poly14_shifted[133]) );
  CFD2QXL \Poly14_reg[273]  ( .D(n10132), .CP(clk), .CD(n18397), .Q(
        poly14_shifted[289]) );
  CFD2QXL \Poly14_reg[184]  ( .D(n10221), .CP(clk), .CD(n18397), .Q(
        poly14_shifted[200]) );
  CFD2QXL \Poly7_reg[318]  ( .D(n9786), .CP(clk), .CD(n18397), .Q(
        poly7_shifted[330]) );
  CFD2QXL \Poly7_reg[146]  ( .D(n9958), .CP(clk), .CD(n18397), .Q(
        poly7_shifted[158]) );
  CFD2QXL \Poly7_reg[337]  ( .D(n9767), .CP(clk), .CD(n18397), .Q(
        poly7_shifted[349]) );
  CFD2QXL \Poly15_reg[0]  ( .D(n9637), .CP(clk), .CD(n18396), .Q(
        poly15_shifted[15]) );
  CFD2QXL \Poly15_reg[7]  ( .D(n9630), .CP(clk), .CD(n18396), .Q(
        poly15_shifted[22]) );
  CFD2QXL \Poly1_reg[302]  ( .D(n9055), .CP(clk), .CD(n18392), .Q(
        poly1_shifted[313]) );
  CFD2QXL \Poly2_reg[4]  ( .D(n9006), .CP(clk), .CD(n18391), .Q(
        poly2_shifted[16]) );
  CFD2QXL \Poly3_reg[6]  ( .D(n8934), .CP(clk), .CD(n18390), .Q(
        poly3_shifted[20]) );
  CFD2QXL \Poly3_reg[8]  ( .D(n8932), .CP(clk), .CD(n18390), .Q(
        poly3_shifted[22]) );
  CFD2QXL \Poly4_reg[11]  ( .D(n8845), .CP(clk), .CD(n18256), .Q(
        poly4_shifted[28]) );
  CFD2QXL \scrambler_reg[4]  ( .D(n8704), .CP(clk), .CD(n18401), .Q(
        scrambler[4]) );
  CFD2QXL \Poly12_reg[4]  ( .D(n10528), .CP(clk), .CD(n18294), .Q(
        poly12_shifted[20]) );
  CFD2QXL \Poly2_reg[44]  ( .D(n8966), .CP(clk), .CD(n18390), .Q(
        poly2_shifted[56]) );
  CFD2QXL \Poly12_reg[73]  ( .D(n10459), .CP(clk), .CD(n18398), .Q(
        poly12_shifted[89]) );
  CFD2QXL \Poly1_reg[300]  ( .D(n9057), .CP(clk), .CD(n18369), .Q(
        poly1_shifted[311]) );
  CFD2QXL \Poly13_reg[493]  ( .D(n10567), .CP(clk), .CD(n18284), .Q(
        poly13_shifted[507]) );
  CFD2QXL \Poly4_reg[33]  ( .D(n8823), .CP(clk), .CD(n18256), .Q(Poly4[33]) );
  CFD2QXL \Poly1_reg[236]  ( .D(n9121), .CP(clk), .CD(n18254), .Q(
        poly1_shifted[247]) );
  CFD2QXL \Poly4_reg[4]  ( .D(n8852), .CP(clk), .CD(n18389), .Q(
        poly4_shifted[21]) );
  CFD2QXL \Poly5_reg[86]  ( .D(n11440), .CP(clk), .CD(n18258), .Q(Poly5[86])
         );
  CFD2QXL \Poly5_reg[80]  ( .D(n11446), .CP(clk), .CD(n18260), .Q(Poly5[80])
         );
  CFD2QXL \Poly12_reg[16]  ( .D(n10516), .CP(clk), .CD(n18292), .Q(Poly12[16])
         );
  CFD2QXL \Poly6_reg[27]  ( .D(n9666), .CP(clk), .CD(n18343), .Q(Poly6[27]) );
  CFD2QXL \Poly2_reg[37]  ( .D(n8973), .CP(clk), .CD(n18391), .Q(Poly2[37]) );
  CFD2QXL \Poly4_reg[25]  ( .D(n8831), .CP(clk), .CD(n18256), .Q(Poly4[25]) );
  CFD2QXL \Poly3_reg[81]  ( .D(n8859), .CP(clk), .CD(n18384), .Q(Poly3[81]) );
  CFD2QXL \Poly14_reg[162]  ( .D(n10243), .CP(clk), .CD(n18398), .Q(
        poly14_shifted[178]) );
  CFD2QXL \Poly1_reg[120]  ( .D(n9237), .CP(clk), .CD(n18392), .Q(
        poly1_shifted[131]) );
  CFD2QXL \Poly1_reg[116]  ( .D(n9241), .CP(clk), .CD(n18392), .Q(
        poly1_shifted[127]) );
  CFD2QXL \Poly3_reg[13]  ( .D(n8927), .CP(clk), .CD(n18390), .Q(
        poly3_shifted[27]) );
  CFD2QXL \Poly1_reg[56]  ( .D(n9301), .CP(clk), .CD(n18392), .Q(Poly1[56]) );
  CFD2QXL \Poly5_reg[121]  ( .D(n11405), .CP(clk), .CD(n18260), .Q(Poly5[121])
         );
  CFD2QXL \Poly2_reg[5]  ( .D(n9005), .CP(clk), .CD(n18391), .Q(
        poly2_shifted[17]) );
  CFD2QXL \Poly11_reg[54]  ( .D(n11135), .CP(clk), .CD(n18257), .Q(Poly11[54])
         );
  CFD2QXL \Poly15_reg[14]  ( .D(n9623), .CP(clk), .CD(n18345), .Q(Poly15[14])
         );
  CFD2QXL \Poly15_reg[13]  ( .D(n9624), .CP(clk), .CD(n18256), .Q(Poly15[13])
         );
  CFD2QXL \Poly11_reg[36]  ( .D(n11153), .CP(clk), .CD(n18257), .Q(Poly11[36])
         );
  CFD2QXL \Poly11_reg[53]  ( .D(n11136), .CP(clk), .CD(n18257), .Q(Poly11[53])
         );
  CFD2QXL \Poly8_reg[8]  ( .D(n11393), .CP(clk), .CD(n18261), .Q(Poly8[8]) );
  CFD2QXL \Poly6_reg[28]  ( .D(n9665), .CP(clk), .CD(n18396), .Q(Poly6[28]) );
  CFD2QXL \Poly0_reg[116]  ( .D(n9461), .CP(clk), .CD(n18350), .Q(Poly0[116])
         );
  CFD2QXL \Poly4_reg[21]  ( .D(n8835), .CP(clk), .CD(n18385), .Q(Poly4[21]) );
  CFD2QXL \Poly12_reg[106]  ( .D(n10426), .CP(clk), .CD(n18293), .Q(
        poly12_shifted[122]) );
  CFD2QXL \Poly12_reg[8]  ( .D(n10524), .CP(clk), .CD(n18398), .Q(
        poly12_shifted[24]) );
  CFD2QXL \Poly3_reg[9]  ( .D(n8931), .CP(clk), .CD(n18390), .Q(
        poly3_shifted[23]) );
  CFD2QXL \Poly3_reg[1]  ( .D(n8939), .CP(clk), .CD(n18390), .Q(
        poly3_shifted[15]) );
  CFD2QXL \dataselector_reg[56]  ( .D(n8739), .CP(clk), .CD(n18402), .Q(
        dataselector[56]) );
  CFD2QXL \dataselector_reg[44]  ( .D(n8751), .CP(clk), .CD(n18257), .Q(
        dataselector[44]) );
  CFD2QXL \Poly12_reg[43]  ( .D(n10489), .CP(clk), .CD(n18296), .Q(
        poly12_shifted[59]) );
  CFD2QXL \Poly3_reg[58]  ( .D(n8882), .CP(clk), .CD(n18390), .Q(Poly3[58]) );
  CFD2QXL \Poly2_reg[30]  ( .D(n8980), .CP(clk), .CD(n18391), .Q(Poly2[30]) );
  CFD2QXL \Poly3_reg[53]  ( .D(n8887), .CP(clk), .CD(n18390), .Q(Poly3[53]) );
  CFD2QXL \Poly4_reg[37]  ( .D(n8819), .CP(clk), .CD(n18389), .Q(Poly4[37]) );
  CFD2QXL \Poly4_reg[35]  ( .D(n8821), .CP(clk), .CD(n18389), .Q(Poly4[35]) );
  CFD2QXL \Poly8_reg[54]  ( .D(n11347), .CP(clk), .CD(n18261), .Q(
        poly8_shifted[68]) );
  CFD2QXL \Poly8_reg[52]  ( .D(n11349), .CP(clk), .CD(n18257), .Q(
        poly8_shifted[66]) );
  CFD2QXL \Poly8_reg[61]  ( .D(n11340), .CP(clk), .CD(n18257), .Q(
        poly8_shifted[75]) );
  CFD2QXL \Poly8_reg[45]  ( .D(n11356), .CP(clk), .CD(n18257), .Q(
        poly8_shifted[59]) );
  CFD2QXL \Poly9_reg[65]  ( .D(n11240), .CP(clk), .CD(n18257), .Q(
        poly9_shifted[76]) );
  CFD2QXL \Poly9_reg[76]  ( .D(n11229), .CP(clk), .CD(n18257), .Q(
        poly9_shifted[87]) );
  CFD2QXL \Poly9_reg[57]  ( .D(n11248), .CP(clk), .CD(n18257), .Q(
        poly9_shifted[68]) );
  CFD2QXL \Poly9_reg[40]  ( .D(n11265), .CP(clk), .CD(n18257), .Q(
        poly9_shifted[51]) );
  CFD2QXL \Poly9_reg[37]  ( .D(n11268), .CP(clk), .CD(n18257), .Q(
        poly9_shifted[48]) );
  CFD2QXL \Poly13_reg[266]  ( .D(n10794), .CP(clk), .CD(n18265), .Q(
        poly13_shifted[280]) );
  CFD2QXL \Poly13_reg[212]  ( .D(n10848), .CP(clk), .CD(n18271), .Q(
        poly13_shifted[226]) );
  CFD2QXL \Poly13_reg[443]  ( .D(n10617), .CP(clk), .CD(n18274), .Q(
        poly13_shifted[457]) );
  CFD2QXL \Poly13_reg[174]  ( .D(n10886), .CP(clk), .CD(n18290), .Q(
        poly13_shifted[188]) );
  CFD2QXL \Poly12_reg[3]  ( .D(n10529), .CP(clk), .CD(n18293), .Q(
        poly12_shifted[19]) );
  CFD2QXL \Poly12_reg[68]  ( .D(n10464), .CP(clk), .CD(n18298), .Q(
        poly12_shifted[84]) );
  CFD2QXL \Poly14_reg[139]  ( .D(n10266), .CP(clk), .CD(n18304), .Q(
        poly14_shifted[155]) );
  CFD2QXL \Poly14_reg[237]  ( .D(n10168), .CP(clk), .CD(n18310), .Q(
        poly14_shifted[253]) );
  CFD2QXL \Poly14_reg[231]  ( .D(n10174), .CP(clk), .CD(n18310), .Q(
        poly14_shifted[247]) );
  CFD2QXL \Poly14_reg[154]  ( .D(n10251), .CP(clk), .CD(n18311), .Q(
        poly14_shifted[170]) );
  CFD2QXL \Poly7_reg[320]  ( .D(n9784), .CP(clk), .CD(n18322), .Q(
        poly7_shifted[332]) );
  CFD2QXL \Poly7_reg[310]  ( .D(n9794), .CP(clk), .CD(n18323), .Q(
        poly7_shifted[322]) );
  CFD2QXL \Poly7_reg[47]  ( .D(n10057), .CP(clk), .CD(n18328), .Q(
        poly7_shifted[59]) );
  CFD2QXL \Poly7_reg[222]  ( .D(n9882), .CP(clk), .CD(n18335), .Q(
        poly7_shifted[234]) );
  CFD2QXL \Poly7_reg[118]  ( .D(n9986), .CP(clk), .CD(n18338), .Q(
        poly7_shifted[130]) );
  CFD2QXL \Poly7_reg[267]  ( .D(n9837), .CP(clk), .CD(n18339), .Q(
        poly7_shifted[279]) );
  CFD2QXL \Poly6_reg[45]  ( .D(n9648), .CP(clk), .CD(n18342), .Q(
        poly6_shifted[55]) );
  CFD2QXL \Poly15_reg[8]  ( .D(n9629), .CP(clk), .CD(n18345), .Q(
        poly15_shifted[23]) );
  CFD2QXL \Poly15_reg[37]  ( .D(n9600), .CP(clk), .CD(n18346), .Q(
        poly15_shifted[52]) );
  CFD2QXL \Poly15_reg[5]  ( .D(n9632), .CP(clk), .CD(n18346), .Q(
        poly15_shifted[20]) );
  CFD2QXL \Poly0_reg[123]  ( .D(n9454), .CP(clk), .CD(n18355), .Q(
        poly0_shifted[141]) );
  CFD2QXL \Poly1_reg[319]  ( .D(n9038), .CP(clk), .CD(n18360), .Q(
        poly1_shifted[330]) );
  CFD2QXL \Poly1_reg[307]  ( .D(n9050), .CP(clk), .CD(n18360), .Q(
        poly1_shifted[318]) );
  CFD2QXL \Poly1_reg[284]  ( .D(n9073), .CP(clk), .CD(n18361), .Q(
        poly1_shifted[295]) );
  CFD2QXL \Poly1_reg[295]  ( .D(n9062), .CP(clk), .CD(n18361), .Q(
        poly1_shifted[306]) );
  CFD2QXL \Poly1_reg[222]  ( .D(n9135), .CP(clk), .CD(n18364), .Q(
        poly1_shifted[233]) );
  CFD2QXL \Poly1_reg[304]  ( .D(n9053), .CP(clk), .CD(n18364), .Q(
        poly1_shifted[315]) );
  CFD2QXL \Poly2_reg[8]  ( .D(n9002), .CP(clk), .CD(n18378), .Q(
        poly2_shifted[20]) );
  CFD2QXL \Poly3_reg[3]  ( .D(n8937), .CP(clk), .CD(n18380), .Q(
        poly3_shifted[17]) );
  CFD2QXL \Poly3_reg[30]  ( .D(n8910), .CP(clk), .CD(n18383), .Q(
        poly3_shifted[44]) );
  CFD2QXL \Poly11_reg[48]  ( .D(n11141), .CP(clk), .CD(n18257), .Q(Poly11[48])
         );
  CFD2QXL \Poly8_reg[22]  ( .D(n11379), .CP(clk), .CD(n18257), .Q(
        poly8_shifted[36]) );
  CFD2QXL \Poly8_reg[64]  ( .D(n11337), .CP(clk), .CD(n18257), .Q(
        poly8_shifted[78]) );
  CFD2QXL \Poly8_reg[21]  ( .D(n11380), .CP(clk), .CD(n18257), .Q(
        poly8_shifted[35]) );
  CFD2QXL \Poly8_reg[63]  ( .D(n11338), .CP(clk), .CD(n18257), .Q(
        poly8_shifted[77]) );
  CFD2QXL \Poly9_reg[11]  ( .D(n11294), .CP(clk), .CD(n18257), .Q(
        poly9_shifted[22]) );
  CFD2QXL \Poly9_reg[101]  ( .D(n11204), .CP(clk), .CD(n18257), .Q(
        poly9_shifted[112]) );
  CFD2QXL \Poly9_reg[69]  ( .D(n11236), .CP(clk), .CD(n18257), .Q(
        poly9_shifted[80]) );
  CFD2QXL \Poly9_reg[80]  ( .D(n11225), .CP(clk), .CD(n18257), .Q(
        poly9_shifted[91]) );
  CFD2QXL \Poly11_reg[0]  ( .D(n11189), .CP(clk), .CD(n18257), .Q(
        poly11_shifted[15]) );
  CFD2QXL \Poly13_reg[487]  ( .D(n10573), .CP(clk), .CD(n18270), .Q(
        poly13_shifted[501]) );
  CFD2QXL \Poly13_reg[268]  ( .D(n10792), .CP(clk), .CD(n18271), .Q(
        poly13_shifted[282]) );
  CFD2QXL \Poly13_reg[206]  ( .D(n10854), .CP(clk), .CD(n18282), .Q(
        poly13_shifted[220]) );
  CFD2QXL \Poly13_reg[376]  ( .D(n10684), .CP(clk), .CD(n18283), .Q(
        poly13_shifted[390]) );
  CFD2QXL \Poly13_reg[219]  ( .D(n10841), .CP(clk), .CD(n18255), .Q(
        poly13_shifted[233]) );
  CFD2QXL \Poly13_reg[506]  ( .D(n10554), .CP(clk), .CD(n18287), .Q(
        poly13_shifted[520]) );
  CFD2QXL \Poly14_reg[61]  ( .D(n10344), .CP(clk), .CD(n18301), .Q(
        poly14_shifted[77]) );
  CFD2QXL \Poly14_reg[75]  ( .D(n10330), .CP(clk), .CD(n18304), .Q(
        poly14_shifted[91]) );
  CFD2QXL \Poly14_reg[281]  ( .D(n10124), .CP(clk), .CD(n18307), .Q(
        poly14_shifted[297]) );
  CFD2QXL \Poly14_reg[253]  ( .D(n10152), .CP(clk), .CD(n18310), .Q(
        poly14_shifted[269]) );
  CFD2QXL \Poly14_reg[50]  ( .D(n10355), .CP(clk), .CD(n18315), .Q(
        poly14_shifted[66]) );
  CFD2QXL \Poly7_reg[398]  ( .D(n9706), .CP(clk), .CD(n18319), .Q(
        poly7_shifted[410]) );
  CFD2QXL \Poly7_reg[368]  ( .D(n9736), .CP(clk), .CD(n18322), .Q(
        poly7_shifted[380]) );
  CFD2QXL \Poly7_reg[307]  ( .D(n9797), .CP(clk), .CD(n18327), .Q(
        poly7_shifted[319]) );
  CFD2QXL \Poly7_reg[140]  ( .D(n9964), .CP(clk), .CD(n18335), .Q(
        poly7_shifted[152]) );
  CFD2QXL \Poly15_reg[40]  ( .D(n9597), .CP(clk), .CD(n18256), .Q(
        poly15_shifted[55]) );
  CFD2QXL \Poly1_reg[264]  ( .D(n9093), .CP(clk), .CD(n18359), .Q(
        poly1_shifted[275]) );
  CFD2QXL \Poly1_reg[90]  ( .D(n9267), .CP(clk), .CD(n18363), .Q(
        poly1_shifted[101]) );
  CFD2QXL \Poly1_reg[249]  ( .D(n9108), .CP(clk), .CD(n18364), .Q(
        poly1_shifted[260]) );
  CFD2QXL \Poly1_reg[89]  ( .D(n9268), .CP(clk), .CD(n18365), .Q(
        poly1_shifted[100]) );
  CFD2QXL \Poly1_reg[248]  ( .D(n9109), .CP(clk), .CD(n18254), .Q(
        poly1_shifted[259]) );
  CFD2QXL \Poly2_reg[1]  ( .D(n9009), .CP(clk), .CD(n18391), .Q(
        poly2_shifted[13]) );
  CFD2QXL \Poly3_reg[25]  ( .D(n8915), .CP(clk), .CD(n18384), .Q(
        poly3_shifted[39]) );
  CFD2QXL \dataselector_reg[40]  ( .D(n8755), .CP(clk), .CD(n18402), .Q(
        dataselector[40]) );
  CFD2QXL \Poly5_reg[116]  ( .D(n11410), .CP(clk), .CD(n18258), .Q(Poly5[116])
         );
  CFD2QXL \Poly13_reg[168]  ( .D(n10892), .CP(clk), .CD(n18265), .Q(
        Poly13[168]) );
  CFD2QXL \Poly5_reg[120]  ( .D(n11406), .CP(clk), .CD(n18258), .Q(Poly5[120])
         );
  CFD2QXL \Poly8_reg[41]  ( .D(n11360), .CP(clk), .CD(n18261), .Q(
        poly8_shifted[55]) );
  CFD2QXL \Poly8_reg[59]  ( .D(n11342), .CP(clk), .CD(n18257), .Q(
        poly8_shifted[73]) );
  CFD2QXL \Poly13_reg[67]  ( .D(n10993), .CP(clk), .CD(n18277), .Q(
        poly13_shifted[81]) );
  CFD2QXL \Poly14_reg[52]  ( .D(n10353), .CP(clk), .CD(n18312), .Q(
        poly14_shifted[68]) );
  CFD2QXL \Poly7_reg[134]  ( .D(n9970), .CP(clk), .CD(n18326), .Q(
        poly7_shifted[146]) );
  CFD2QXL \scrambler_reg[6]  ( .D(n8706), .CP(clk), .CD(n18401), .Q(
        scrambler[6]) );
  CFD2QXL \scrambler_reg[3]  ( .D(n8703), .CP(clk), .CD(n18257), .Q(
        scrambler[3]) );
  CFD2QXL \scrambler_reg[0]  ( .D(n8700), .CP(clk), .CD(n18401), .Q(
        scrambler[0]) );
  CFD2QXL \Poly11_reg[21]  ( .D(n11168), .CP(clk), .CD(n18257), .Q(Poly11[21])
         );
  CFD2QXL \Poly3_reg[65]  ( .D(n8875), .CP(clk), .CD(n18381), .Q(
        poly3_shifted[79]) );
  CFD2QXL \Poly11_reg[11]  ( .D(n11178), .CP(clk), .CD(n18257), .Q(
        poly11_shifted[26]) );
  CFD2QXL \Poly6_reg[50]  ( .D(n9643), .CP(clk), .CD(n18341), .Q(Poly6[50]) );
  CFD2QXL \Poly2_reg[11]  ( .D(n8999), .CP(clk), .CD(n18378), .Q(
        poly2_shifted[23]) );
  CFD2QXL \Poly13_reg[385]  ( .D(n10675), .CP(clk), .CD(n18288), .Q(
        poly13_shifted[399]) );
  CFD2QXL \Poly0_reg[125]  ( .D(n9452), .CP(clk), .CD(n18356), .Q(
        poly0_shifted[143]) );
  CFD2QXL \Poly1_reg[103]  ( .D(n9254), .CP(clk), .CD(n18376), .Q(
        poly1_shifted[114]) );
  CFD2QXL \Poly9_reg[48]  ( .D(n11257), .CP(clk), .CD(n18257), .Q(
        poly9_shifted[59]) );
  CFD2QXL \scrambler_reg[13]  ( .D(n8713), .CP(clk), .CD(n18257), .Q(
        scrambler[13]) );
  CFD2QXL \scrambler_reg[2]  ( .D(n8702), .CP(clk), .CD(n18401), .Q(
        scrambler[2]) );
  CFD2QXL \Poly0_reg[211]  ( .D(n9366), .CP(clk), .CD(n18352), .Q(Poly0[211])
         );
  CFD2QXL \Poly8_reg[2]  ( .D(n11399), .CP(clk), .CD(n18257), .Q(Poly8[2]) );
  CFD2QXL \Poly12_reg[95]  ( .D(n10437), .CP(clk), .CD(n18298), .Q(Poly12[95])
         );
  CFD2QXL \Poly7_reg[178]  ( .D(n9926), .CP(clk), .CD(n18338), .Q(Poly7[178])
         );
  CFD2QXL \Poly3_reg[31]  ( .D(n8909), .CP(clk), .CD(n18380), .Q(Poly3[31]) );
  CFD2QXL \Poly4_reg[16]  ( .D(n8840), .CP(clk), .CD(n18384), .Q(Poly4[16]) );
  CFD2QXL \dataselector_reg[37]  ( .D(n8758), .CP(clk), .CD(n18257), .Q(
        dataselector[37]) );
  CFD2QXL \scrambler_reg[7]  ( .D(n8707), .CP(clk), .CD(n18257), .Q(
        scrambler[7]) );
  CFD2QXL \Poly8_reg[68]  ( .D(n11333), .CP(clk), .CD(n18261), .Q(Poly8[68])
         );
  CFD2QXL \Poly8_reg[76]  ( .D(n11325), .CP(clk), .CD(n18257), .Q(Poly8[76])
         );
  CFD2QXL \Poly7_reg[25]  ( .D(n10079), .CP(clk), .CD(n18320), .Q(Poly7[25])
         );
  CFD2QXL \Poly4_reg[26]  ( .D(n8830), .CP(clk), .CD(n18385), .Q(Poly4[26]) );
  CFD2QXL \Poly0_reg[110]  ( .D(n9467), .CP(clk), .CD(n18355), .Q(Poly0[110])
         );
  CFD2QXL \Poly2_reg[42]  ( .D(n8968), .CP(clk), .CD(n18379), .Q(Poly2[42]) );
  CFD2QXL \Poly9_reg[24]  ( .D(n11281), .CP(clk), .CD(n18257), .Q(Poly9[24])
         );
  CFD2QXL \Poly11_reg[43]  ( .D(n11146), .CP(clk), .CD(n18257), .Q(Poly11[43])
         );
  CFD2QXL \Poly6_reg[4]  ( .D(n9689), .CP(clk), .CD(n18342), .Q(Poly6[4]) );
  CFD2QXL \Poly2_reg[41]  ( .D(n8969), .CP(clk), .CD(n18391), .Q(Poly2[41]) );
  CFD2QXL \Poly6_reg[43]  ( .D(n9650), .CP(clk), .CD(n18344), .Q(Poly6[43]) );
  CFD2QXL \Poly10_reg[14]  ( .D(n11089), .CP(clk), .CD(n18263), .Q(Poly10[14])
         );
  CFD2QXL \Poly6_reg[18]  ( .D(n9675), .CP(clk), .CD(n18342), .Q(Poly6[18]) );
  CFD2QXL \Poly10_reg[36]  ( .D(n11067), .CP(clk), .CD(n18262), .Q(Poly10[36])
         );
  CFD2QXL \Poly14_reg[177]  ( .D(n10228), .CP(clk), .CD(n18303), .Q(
        Poly14[177]) );
  CFD2QXL \Poly6_reg[51]  ( .D(n9642), .CP(clk), .CD(n18344), .Q(Poly6[51]) );
  CFD2QXL \Poly6_reg[54]  ( .D(n9639), .CP(clk), .CD(n18342), .Q(Poly6[54]) );
  CFD2QXL \Poly6_reg[7]  ( .D(n9686), .CP(clk), .CD(n18343), .Q(
        poly6_shifted[17]) );
  CFD2QXL \Poly2_reg[25]  ( .D(n8985), .CP(clk), .CD(n18379), .Q(Poly2[25]) );
  CFD2QXL \Poly6_reg[14]  ( .D(n9679), .CP(clk), .CD(n18342), .Q(Poly6[14]) );
  CFD2QXL \Poly0_reg[197]  ( .D(n9380), .CP(clk), .CD(n18354), .Q(
        poly0_shifted[215]) );
  CFD2QXL \Poly15_reg[28]  ( .D(n9609), .CP(clk), .CD(n18256), .Q(Poly15[28])
         );
  CFD2QXL \Poly0_reg[199]  ( .D(n9378), .CP(clk), .CD(n18355), .Q(
        poly0_shifted[217]) );
  CFD2QXL \Poly15_reg[27]  ( .D(n9610), .CP(clk), .CD(n18345), .Q(Poly15[27])
         );
  CFD2QXL \Poly15_reg[16]  ( .D(n9621), .CP(clk), .CD(n18345), .Q(Poly15[16])
         );
  CFD2QXL \Poly5_reg[122]  ( .D(n11404), .CP(clk), .CD(n18257), .Q(Poly5[122])
         );
  CFD2QXL \Poly0_reg[212]  ( .D(n9365), .CP(clk), .CD(n18349), .Q(Poly0[212])
         );
  CFD2QXL \Poly6_reg[26]  ( .D(n9667), .CP(clk), .CD(n18344), .Q(Poly6[26]) );
  CFD2QXL \Poly11_reg[73]  ( .D(n11116), .CP(clk), .CD(n18257), .Q(Poly11[73])
         );
  CFD2QXL \Poly6_reg[25]  ( .D(n9668), .CP(clk), .CD(n18344), .Q(Poly6[25]) );
  CFD2QXL \Poly10_reg[0]  ( .D(n11103), .CP(clk), .CD(n18400), .Q(Poly10[0])
         );
  CFD2QXL \Poly10_reg[22]  ( .D(n11081), .CP(clk), .CD(n18263), .Q(Poly10[22])
         );
  CFD2QXL \Poly9_reg[44]  ( .D(n11261), .CP(clk), .CD(n18257), .Q(
        poly9_shifted[55]) );
  CFD2QXL \Poly12_reg[89]  ( .D(n10443), .CP(clk), .CD(n18398), .Q(Poly12[89])
         );
  CFD2QXL \Poly7_reg[378]  ( .D(n9726), .CP(clk), .CD(n18397), .Q(
        poly7_shifted[390]) );
  CFD2QXL \Poly6_reg[30]  ( .D(n9663), .CP(clk), .CD(n18341), .Q(Poly6[30]) );
  CFD2QXL \Poly1_reg[154]  ( .D(n9203), .CP(clk), .CD(n18392), .Q(Poly1[154])
         );
  CFD2QXL \Poly1_reg[228]  ( .D(n9129), .CP(clk), .CD(n18392), .Q(Poly1[228])
         );
  CFD2QXL \Poly1_reg[201]  ( .D(n9156), .CP(clk), .CD(n18392), .Q(Poly1[201])
         );
  CFD2QXL \Poly6_reg[1]  ( .D(n9692), .CP(clk), .CD(n18342), .Q(Poly6[1]) );
  CFD2QXL \Poly6_reg[11]  ( .D(n9682), .CP(clk), .CD(n18343), .Q(Poly6[11]) );
  CFD2QXL \Poly2_reg[56]  ( .D(n8954), .CP(clk), .CD(n18390), .Q(Poly2[56]) );
  CFD2QXL \Poly6_reg[33]  ( .D(n9660), .CP(clk), .CD(n18344), .Q(Poly6[33]) );
  CFD2QXL \Poly11_reg[71]  ( .D(n11118), .CP(clk), .CD(n18257), .Q(Poly11[71])
         );
  CFD2QXL \Poly5_reg[36]  ( .D(n11490), .CP(clk), .CD(n18259), .Q(
        poly5_shifted[50]) );
  CFD2QXL \Poly15_reg[59]  ( .D(n9578), .CP(clk), .CD(n18396), .Q(Poly15[59])
         );
  CFD2QXL \Poly1_reg[339]  ( .D(n9018), .CP(clk), .CD(n18393), .Q(Poly1[339])
         );
  CFD2QXL \Poly3_reg[39]  ( .D(n8901), .CP(clk), .CD(n18384), .Q(Poly3[39]) );
  CFD2QXL \Poly0_reg[11]  ( .D(n9566), .CP(clk), .CD(n18396), .Q(Poly0[11]) );
  CFD2QXL \Poly1_reg[149]  ( .D(n9208), .CP(clk), .CD(n18392), .Q(
        poly1_shifted[160]) );
  CFD2QXL \Poly7_reg[212]  ( .D(n9892), .CP(clk), .CD(n18397), .Q(
        poly7_shifted[224]) );
  CFD2QXL \Poly5_reg[85]  ( .D(n11441), .CP(clk), .CD(n18257), .Q(Poly5[85])
         );
  CFD2QXL \Poly3_reg[7]  ( .D(n8933), .CP(clk), .CD(n18382), .Q(
        poly3_shifted[21]) );
  CFD2QXL \Poly9_reg[56]  ( .D(n11249), .CP(clk), .CD(n18257), .Q(
        poly9_shifted[67]) );
  CFD2QXL \Poly13_reg[119]  ( .D(n10941), .CP(clk), .CD(n18399), .Q(
        poly13_shifted[133]) );
  CFD2QXL \Poly15_reg[9]  ( .D(n9628), .CP(clk), .CD(n18346), .Q(
        poly15_shifted[24]) );
  CFD2QXL \Poly2_reg[62]  ( .D(n8948), .CP(clk), .CD(n18392), .Q(Poly2[62]) );
  CFD2QXL \Poly11_reg[32]  ( .D(n11157), .CP(clk), .CD(n18257), .Q(Poly11[32])
         );
  CFD2QXL \Poly11_reg[35]  ( .D(n11154), .CP(clk), .CD(n18257), .Q(Poly11[35])
         );
  CFD2QXL \Poly10_reg[37]  ( .D(n11066), .CP(clk), .CD(n18263), .Q(Poly10[37])
         );
  CFD2QXL \Poly8_reg[82]  ( .D(n11319), .CP(clk), .CD(n18257), .Q(Poly8[82])
         );
  CFD2QXL \Poly8_reg[67]  ( .D(n11334), .CP(clk), .CD(n18257), .Q(Poly8[67])
         );
  CFD2QXL \Poly14_reg[198]  ( .D(n10207), .CP(clk), .CD(n18309), .Q(
        Poly14[198]) );
  CFD2QXL \Poly1_reg[61]  ( .D(n9296), .CP(clk), .CD(n18375), .Q(Poly1[61]) );
  CFD2QXL \Poly15_reg[33]  ( .D(n9604), .CP(clk), .CD(n18396), .Q(Poly15[33])
         );
  CFD2QXL \Poly12_reg[91]  ( .D(n10441), .CP(clk), .CD(n18297), .Q(Poly12[91])
         );
  CFD2QXL \Poly6_reg[20]  ( .D(n9673), .CP(clk), .CD(n18341), .Q(Poly6[20]) );
  CFD2QXL \Poly6_reg[42]  ( .D(n9651), .CP(clk), .CD(n18343), .Q(Poly6[42]) );
  CFD2QXL \Poly6_reg[24]  ( .D(n9669), .CP(clk), .CD(n18396), .Q(Poly6[24]) );
  CFD2QXL \Poly15_reg[31]  ( .D(n9606), .CP(clk), .CD(n18396), .Q(Poly15[31])
         );
  CFD2QXL \Poly2_reg[38]  ( .D(n8972), .CP(clk), .CD(n18391), .Q(Poly2[38]) );
  CFD2QXL \Poly2_reg[60]  ( .D(n8950), .CP(clk), .CD(n18391), .Q(Poly2[60]) );
  CFD2QXL \Poly2_reg[58]  ( .D(n8952), .CP(clk), .CD(n18391), .Q(Poly2[58]) );
  CFD2QXL \Poly11_reg[67]  ( .D(n11122), .CP(clk), .CD(n18257), .Q(Poly11[67])
         );
  CFD2QXL \Poly8_reg[73]  ( .D(n11328), .CP(clk), .CD(n18257), .Q(Poly8[73])
         );
  CFD2QXL \Poly11_reg[72]  ( .D(n11117), .CP(clk), .CD(n18262), .Q(Poly11[72])
         );
  CFD2QXL \Poly12_reg[112]  ( .D(n10420), .CP(clk), .CD(n18292), .Q(
        Poly12[112]) );
  CFD2QXL \Poly11_reg[40]  ( .D(n11149), .CP(clk), .CD(n18257), .Q(Poly11[40])
         );
  CFD2QXL \Poly6_reg[46]  ( .D(n9647), .CP(clk), .CD(n18397), .Q(Poly6[46]) );
  CFD2QXL \Poly12_reg[111]  ( .D(n10421), .CP(clk), .CD(n18297), .Q(
        Poly12[111]) );
  CFD2QXL \Poly12_reg[122]  ( .D(n10410), .CP(clk), .CD(n18293), .Q(
        Poly12[122]) );
  CFD2QXL \Poly12_reg[124]  ( .D(n10408), .CP(clk), .CD(n18294), .Q(
        Poly12[124]) );
  CFD2QXL \Poly6_reg[47]  ( .D(n9646), .CP(clk), .CD(n18342), .Q(Poly6[47]) );
  CFD2QXL \Poly10_reg[34]  ( .D(n11069), .CP(clk), .CD(n18263), .Q(Poly10[34])
         );
  CFD2QXL \Poly7_reg[399]  ( .D(n9705), .CP(clk), .CD(n18339), .Q(Poly7[399])
         );
  CFD2QXL \Poly10_reg[25]  ( .D(n11078), .CP(clk), .CD(n18263), .Q(Poly10[25])
         );
  CFD2QXL \Poly2_reg[63]  ( .D(n8947), .CP(clk), .CD(n18392), .Q(Poly2[63]) );
  CFD2QXL \Poly7_reg[404]  ( .D(n9700), .CP(clk), .CD(n18322), .Q(
        \dataselector_shifted[0] ) );
  CFD2QXL \Poly15_reg[32]  ( .D(n9605), .CP(clk), .CD(n18256), .Q(Poly15[32])
         );
  CFD2QXL \Poly0_reg[156]  ( .D(n9421), .CP(clk), .CD(n18394), .Q(Poly0[156])
         );
  CFD2QXL \Poly3_reg[57]  ( .D(n8883), .CP(clk), .CD(n18382), .Q(Poly3[57]) );
  CFD2QXL \Poly12_reg[115]  ( .D(n10417), .CP(clk), .CD(n18294), .Q(
        Poly12[115]) );
  CFD2QXL \Poly1_reg[346]  ( .D(n9011), .CP(clk), .CD(n18393), .Q(Poly1[346])
         );
  CFD2QXL \Poly1_reg[336]  ( .D(n9021), .CP(clk), .CD(n18393), .Q(Poly1[336])
         );
  CFD2QXL \Poly12_reg[116]  ( .D(n10416), .CP(clk), .CD(n18293), .Q(
        Poly12[116]) );
  CFD2QXL \Poly7_reg[403]  ( .D(n9701), .CP(clk), .CD(n18327), .Q(Poly7[403])
         );
  CFD2QXL \Poly12_reg[113]  ( .D(n10419), .CP(clk), .CD(n18399), .Q(
        Poly12[113]) );
  CFD2QXL \Poly8_reg[1]  ( .D(n11400), .CP(clk), .CD(n18257), .Q(Poly8[1]) );
  CFD2QXL \Poly12_reg[31]  ( .D(n10501), .CP(clk), .CD(n18297), .Q(Poly12[31])
         );
  CFD2QXL \Poly6_reg[29]  ( .D(n9664), .CP(clk), .CD(n18342), .Q(Poly6[29]) );
  CFD2QXL \Poly11_reg[39]  ( .D(n11150), .CP(clk), .CD(n18257), .Q(Poly11[39])
         );
  CFD2QXL \Poly6_reg[41]  ( .D(n9652), .CP(clk), .CD(n18344), .Q(Poly6[41]) );
  CFD2QXL \Poly7_reg[402]  ( .D(n9702), .CP(clk), .CD(n18321), .Q(Poly7[402])
         );
  CFD2QXL \Poly7_reg[401]  ( .D(n9703), .CP(clk), .CD(n18325), .Q(Poly7[401])
         );
  CFD2QXL \Poly1_reg[342]  ( .D(n9015), .CP(clk), .CD(n18393), .Q(Poly1[342])
         );
  CFD2QXL \Poly12_reg[123]  ( .D(n10409), .CP(clk), .CD(n18296), .Q(
        Poly12[123]) );
  CFD2QXL \Poly1_reg[340]  ( .D(n9017), .CP(clk), .CD(n18393), .Q(Poly1[340])
         );
  CFD2QXL \Poly1_reg[338]  ( .D(n9019), .CP(clk), .CD(n18393), .Q(Poly1[338])
         );
  CFD2QXL \Poly1_reg[337]  ( .D(n9020), .CP(clk), .CD(n18393), .Q(Poly1[337])
         );
  CFD2QXL \Poly1_reg[343]  ( .D(n9014), .CP(clk), .CD(n18393), .Q(Poly1[343])
         );
  CFD2QXL \Poly12_reg[121]  ( .D(n10411), .CP(clk), .CD(n18295), .Q(
        Poly12[121]) );
  CFD2QXL \Poly12_reg[17]  ( .D(n10515), .CP(clk), .CD(n18398), .Q(Poly12[17])
         );
  CFD2QXL \Poly6_reg[49]  ( .D(n9644), .CP(clk), .CD(n18342), .Q(Poly6[49]) );
  CFD2QXL \Poly7_reg[400]  ( .D(n9704), .CP(clk), .CD(n18320), .Q(Poly7[400])
         );
  CFD2QXL \Poly7_reg[405]  ( .D(n9699), .CP(clk), .CD(n18330), .Q(Poly7[405])
         );
  CFD2QXL \Poly6_reg[53]  ( .D(n9640), .CP(clk), .CD(n18343), .Q(Poly6[53]) );
  CFD2QXL \Poly1_reg[345]  ( .D(n9012), .CP(clk), .CD(n18393), .Q(Poly1[345])
         );
  CFD2QXL \Poly1_reg[344]  ( .D(n9013), .CP(clk), .CD(n18393), .Q(Poly1[344])
         );
  CFD2QXL \Poly10_reg[42]  ( .D(n11061), .CP(clk), .CD(n18264), .Q(Poly10[42])
         );
  CFD2QXL \Poly11_reg[25]  ( .D(n11164), .CP(clk), .CD(n18257), .Q(Poly11[25])
         );
  CFD2QXL \Poly6_reg[16]  ( .D(n9677), .CP(clk), .CD(n18396), .Q(Poly6[16]) );
  CFD2QXL \Poly6_reg[15]  ( .D(n9678), .CP(clk), .CD(n18396), .Q(Poly6[15]) );
  CFD2QXL \Poly3_reg[46]  ( .D(n8894), .CP(clk), .CD(n18382), .Q(Poly3[46]) );
  CFD2QXL \Poly11_reg[49]  ( .D(n11140), .CP(clk), .CD(n18257), .Q(Poly11[49])
         );
  CFD2QXL \Poly11_reg[28]  ( .D(n11161), .CP(clk), .CD(n18257), .Q(Poly11[28])
         );
  CFD2QXL \Poly12_reg[90]  ( .D(n10442), .CP(clk), .CD(n18398), .Q(Poly12[90])
         );
  CFD2QXL \Poly6_reg[0]  ( .D(n9693), .CP(clk), .CD(n18396), .Q(Poly6[0]) );
  CFD2QXL \Poly7_reg[407]  ( .D(n9697), .CP(clk), .CD(n18333), .Q(Poly7[407])
         );
  CFD2QXL \Poly0_reg[109]  ( .D(n9468), .CP(clk), .CD(n18394), .Q(Poly0[109])
         );
  CFD2QXL \Poly7_reg[410]  ( .D(n9694), .CP(clk), .CD(n18319), .Q(Poly7[410])
         );
  CFD2QXL \Poly7_reg[406]  ( .D(n9698), .CP(clk), .CD(n18323), .Q(Poly7[406])
         );
  CFD2QXL \Poly10_reg[39]  ( .D(n11064), .CP(clk), .CD(n18263), .Q(Poly10[39])
         );
  CFD2QXL \Poly15_reg[54]  ( .D(n9583), .CP(clk), .CD(n18396), .Q(Poly15[54])
         );
  CFD2QXL \Poly10_reg[31]  ( .D(n11072), .CP(clk), .CD(n18400), .Q(Poly10[31])
         );
  CFD2QXL \Poly7_reg[408]  ( .D(n9696), .CP(clk), .CD(n18318), .Q(Poly7[408])
         );
  CFD2QXL \Poly3_reg[79]  ( .D(n8861), .CP(clk), .CD(n18381), .Q(Poly3[79]) );
  CFD2QXL \Poly10_reg[40]  ( .D(n11063), .CP(clk), .CD(n18264), .Q(Poly10[40])
         );
  CFD2QXL \Poly7_reg[409]  ( .D(n9695), .CP(clk), .CD(n18336), .Q(Poly7[409])
         );
  CFD2QXL \Poly5_reg[111]  ( .D(n11415), .CP(clk), .CD(n18257), .Q(Poly5[111])
         );
  CFD2QXL \Poly13_reg[519]  ( .D(n10541), .CP(clk), .CD(n18289), .Q(
        Poly13[519]) );
  CFD2QXL \Poly14_reg[296]  ( .D(n10109), .CP(clk), .CD(n18303), .Q(
        Poly14[296]) );
  CFD2QXL \Poly8_reg[87]  ( .D(n11314), .CP(clk), .CD(n18257), .Q(Poly8[87])
         );
  CFD2QXL \Poly8_reg[91]  ( .D(n11310), .CP(clk), .CD(n18261), .Q(Poly8[91])
         );
  CFD2QXL \Poly0_reg[216]  ( .D(n9361), .CP(clk), .CD(n18347), .Q(Poly0[216])
         );
  CFD2QXL \Poly11_reg[61]  ( .D(n11128), .CP(clk), .CD(n18400), .Q(Poly11[61])
         );
  CFD2QXL \Poly14_reg[294]  ( .D(n10111), .CP(clk), .CD(n18306), .Q(
        Poly14[294]) );
  CFD2QXL \Poly12_reg[120]  ( .D(n10412), .CP(clk), .CD(n18399), .Q(
        Poly12[120]) );
  CFD2QXL \Poly8_reg[89]  ( .D(n11312), .CP(clk), .CD(n18261), .Q(Poly8[89])
         );
  CFD2QXL \Poly10_reg[33]  ( .D(n11070), .CP(clk), .CD(n18400), .Q(Poly10[33])
         );
  CFD2QXL \Poly8_reg[92]  ( .D(n11309), .CP(clk), .CD(n18257), .Q(Poly8[92])
         );
  CFD2QXL \Poly13_reg[525]  ( .D(n10535), .CP(clk), .CD(n18277), .Q(
        Poly13[525]) );
  CFD2QXL \Poly3_reg[74]  ( .D(n8866), .CP(clk), .CD(n18382), .Q(Poly3[74]) );
  CFD2QXL \Poly3_reg[83]  ( .D(n8857), .CP(clk), .CD(n18383), .Q(Poly3[83]) );
  CFD2QXL \Poly12_reg[118]  ( .D(n10414), .CP(clk), .CD(n18399), .Q(
        Poly12[118]) );
  CFD2QXL \Poly0_reg[217]  ( .D(n9360), .CP(clk), .CD(n18355), .Q(Poly0[217])
         );
  CFD2QXL \Poly0_reg[203]  ( .D(n9374), .CP(clk), .CD(n18357), .Q(Poly0[203])
         );
  CFD2QXL \Poly0_reg[209]  ( .D(n9368), .CP(clk), .CD(n18351), .Q(Poly0[209])
         );
  CFD2QXL \Poly0_reg[213]  ( .D(n9364), .CP(clk), .CD(n18353), .Q(Poly0[213])
         );
  CFD2QXL \Poly3_reg[76]  ( .D(n8864), .CP(clk), .CD(n18381), .Q(Poly3[76]) );
  CFD2QXL \Poly3_reg[80]  ( .D(n8860), .CP(clk), .CD(n18382), .Q(Poly3[80]) );
  CFD2QXL \Poly3_reg[73]  ( .D(n8867), .CP(clk), .CD(n18380), .Q(Poly3[73]) );
  CFD2QXL \Poly9_reg[111]  ( .D(n11194), .CP(clk), .CD(n18257), .Q(Poly9[111])
         );
  CFD2QXL \Poly15_reg[50]  ( .D(n9587), .CP(clk), .CD(n18346), .Q(Poly15[50])
         );
  CFD2QXL \Poly9_reg[112]  ( .D(n11193), .CP(clk), .CD(n18257), .Q(Poly9[112])
         );
  CFD2QXL \Poly9_reg[113]  ( .D(n11192), .CP(clk), .CD(n18257), .Q(Poly9[113])
         );
  CFD2QXL \Poly15_reg[53]  ( .D(n9584), .CP(clk), .CD(n18345), .Q(Poly15[53])
         );
  CFD2QXL \Poly9_reg[110]  ( .D(n11195), .CP(clk), .CD(n18257), .Q(Poly9[110])
         );
  CFD2QXL \Poly14_reg[291]  ( .D(n10114), .CP(clk), .CD(n18309), .Q(
        Poly14[291]) );
  CFD2QXL \Poly14_reg[293]  ( .D(n10112), .CP(clk), .CD(n18314), .Q(
        Poly14[293]) );
  CFD2QXL \Poly9_reg[115]  ( .D(n11190), .CP(clk), .CD(n18257), .Q(Poly9[115])
         );
  CFD2QXL \Poly0_reg[210]  ( .D(n9367), .CP(clk), .CD(n18348), .Q(Poly0[210])
         );
  CFD2QXL \Poly0_reg[214]  ( .D(n9363), .CP(clk), .CD(n18349), .Q(Poly0[214])
         );
  CFD2QXL \Poly0_reg[205]  ( .D(n9372), .CP(clk), .CD(n18349), .Q(Poly0[205])
         );
  CFD2QXL \Poly0_reg[218]  ( .D(n9359), .CP(clk), .CD(n18347), .Q(Poly0[218])
         );
  CFD2QXL \Poly0_reg[202]  ( .D(n9375), .CP(clk), .CD(n18348), .Q(Poly0[202])
         );
  CFD2QXL \Poly0_reg[215]  ( .D(n9362), .CP(clk), .CD(n18354), .Q(Poly0[215])
         );
  CFD2QXL \Poly15_reg[51]  ( .D(n9586), .CP(clk), .CD(n18256), .Q(Poly15[51])
         );
  CFD2QXL \Poly8_reg[94]  ( .D(n11307), .CP(clk), .CD(n18257), .Q(Poly8[94])
         );
  CFD2QXL \Poly10_reg[41]  ( .D(n11062), .CP(clk), .CD(n18400), .Q(Poly10[41])
         );
  CFD2QXL \Poly8_reg[86]  ( .D(n11315), .CP(clk), .CD(n18257), .Q(Poly8[86])
         );
  CFD2QXL \Poly15_reg[52]  ( .D(n9585), .CP(clk), .CD(n18346), .Q(Poly15[52])
         );
  CFD2QXL \Poly8_reg[84]  ( .D(n11317), .CP(clk), .CD(n18257), .Q(Poly8[84])
         );
  CFD2QXL \Poly2_reg[69]  ( .D(n8941), .CP(clk), .CD(n18378), .Q(Poly2[69]) );
  CFD2QXL \Poly8_reg[95]  ( .D(n11306), .CP(clk), .CD(n18257), .Q(Poly8[95])
         );
  CFD2QXL \Poly14_reg[288]  ( .D(n10117), .CP(clk), .CD(n18254), .Q(
        Poly14[288]) );
  CFD2QXL \Poly8_reg[85]  ( .D(n11316), .CP(clk), .CD(n18257), .Q(Poly8[85])
         );
  CFD2QXL \Poly9_reg[114]  ( .D(n11191), .CP(clk), .CD(n18257), .Q(Poly9[114])
         );
  CFD2QXL \Poly14_reg[289]  ( .D(n10116), .CP(clk), .CD(n18312), .Q(
        Poly14[289]) );
  CFD2QXL \Poly8_reg[93]  ( .D(n11308), .CP(clk), .CD(n18257), .Q(Poly8[93])
         );
  CFD2QXL \Poly14_reg[292]  ( .D(n10113), .CP(clk), .CD(n18301), .Q(
        Poly14[292]) );
  CFD2QXL \Poly8_reg[83]  ( .D(n11318), .CP(clk), .CD(n18257), .Q(Poly8[83])
         );
  CFD2QXL \Poly9_reg[109]  ( .D(n11196), .CP(clk), .CD(n18257), .Q(Poly9[109])
         );
  CFD2QXL \Poly9_reg[108]  ( .D(n11197), .CP(clk), .CD(n18257), .Q(Poly9[108])
         );
  CFD2QXL \Poly14_reg[300]  ( .D(n10105), .CP(clk), .CD(n18305), .Q(
        Poly14[300]) );
  CFD2QXL \Poly15_reg[56]  ( .D(n9581), .CP(clk), .CD(n18346), .Q(Poly15[56])
         );
  CFD2QXL \Poly13_reg[518]  ( .D(n10542), .CP(clk), .CD(n18266), .Q(
        Poly13[518]) );
  CFD2QXL \Poly13_reg[517]  ( .D(n10543), .CP(clk), .CD(n18267), .Q(
        Poly13[517]) );
  CFD2QXL \Poly13_reg[516]  ( .D(n10544), .CP(clk), .CD(n18269), .Q(
        Poly13[516]) );
  CFD2QXL \Poly13_reg[526]  ( .D(n10534), .CP(clk), .CD(n18276), .Q(
        Poly13[526]) );
  CFD2QXL \Poly14_reg[298]  ( .D(n10107), .CP(clk), .CD(n18300), .Q(
        Poly14[298]) );
  CFD2QXL \Poly9_reg[105]  ( .D(n11200), .CP(clk), .CD(n18257), .Q(Poly9[105])
         );
  CFD2QXL \Poly5_reg[124]  ( .D(n11402), .CP(clk), .CD(n18258), .Q(Poly5[124])
         );
  CFD2QXL \Poly3_reg[72]  ( .D(n8868), .CP(clk), .CD(n18383), .Q(Poly3[72]) );
  CFD2QXL \Poly3_reg[75]  ( .D(n8865), .CP(clk), .CD(n18383), .Q(Poly3[75]) );
  CFD2QXL \Poly3_reg[78]  ( .D(n8862), .CP(clk), .CD(n18384), .Q(Poly3[78]) );
  CFD2QXL \Poly0_reg[204]  ( .D(n9373), .CP(clk), .CD(n18348), .Q(Poly0[204])
         );
  CFD2QXL \Poly3_reg[70]  ( .D(n8870), .CP(clk), .CD(n18380), .Q(Poly3[70]) );
  CFD2QXL \Poly14_reg[295]  ( .D(n10110), .CP(clk), .CD(n18310), .Q(
        Poly14[295]) );
  CFD2QXL \Poly5_reg[123]  ( .D(n11403), .CP(clk), .CD(n18257), .Q(Poly5[123])
         );
  CFD2QXL \Poly9_reg[106]  ( .D(n11199), .CP(clk), .CD(n18257), .Q(Poly9[106])
         );
  CFD2QXL \Poly13_reg[514]  ( .D(n10546), .CP(clk), .CD(n18272), .Q(
        Poly13[514]) );
  CFD2QXL \Poly13_reg[523]  ( .D(n10537), .CP(clk), .CD(n18281), .Q(
        Poly13[523]) );
  CFD2QXL \Poly14_reg[299]  ( .D(n10106), .CP(clk), .CD(n18313), .Q(
        Poly14[299]) );
  CFD2QXL \Poly5_reg[118]  ( .D(n11408), .CP(clk), .CD(n18257), .Q(Poly5[118])
         );
  CFD2QXL \Poly13_reg[515]  ( .D(n10545), .CP(clk), .CD(n18270), .Q(
        Poly13[515]) );
  CFD2QXL \Poly5_reg[115]  ( .D(n11411), .CP(clk), .CD(n18257), .Q(Poly5[115])
         );
  CFD2QXL \Poly15_reg[45]  ( .D(n9592), .CP(clk), .CD(n18344), .Q(Poly15[45])
         );
  CFD2QXL \Poly14_reg[286]  ( .D(n10119), .CP(clk), .CD(n18302), .Q(
        Poly14[286]) );
  CFD2QXL \Poly0_reg[207]  ( .D(n9370), .CP(clk), .CD(n18350), .Q(Poly0[207])
         );
  CFD2QXL \Poly3_reg[77]  ( .D(n8863), .CP(clk), .CD(n18390), .Q(Poly3[77]) );
  CFD2QXL \Poly13_reg[522]  ( .D(n10538), .CP(clk), .CD(n18283), .Q(
        Poly13[522]) );
  CFD2QXL \Poly14_reg[290]  ( .D(n10115), .CP(clk), .CD(n18304), .Q(
        Poly14[290]) );
  CFD2QXL \Poly0_reg[219]  ( .D(n9358), .CP(clk), .CD(n18356), .Q(Poly0[219])
         );
  CFD2QXL \Poly15_reg[47]  ( .D(n9590), .CP(clk), .CD(n18256), .Q(Poly15[47])
         );
  CFD2QXL \Poly14_reg[287]  ( .D(n10118), .CP(clk), .CD(n18315), .Q(
        Poly14[287]) );
  CFD2QXL \Poly13_reg[524]  ( .D(n10536), .CP(clk), .CD(n18279), .Q(
        Poly13[524]) );
  CFD2QXL \Poly13_reg[521]  ( .D(n10539), .CP(clk), .CD(n18284), .Q(
        Poly13[521]) );
  CFD2QXL \Poly8_reg[88]  ( .D(n11313), .CP(clk), .CD(n18257), .Q(Poly8[88])
         );
  CFD2QXL \Poly9_reg[107]  ( .D(n11198), .CP(clk), .CD(n18257), .Q(Poly9[107])
         );
  CFD2QXL \Poly14_reg[297]  ( .D(n10108), .CP(clk), .CD(n18307), .Q(
        Poly14[297]) );
  CFD2QXL \Poly15_reg[55]  ( .D(n9582), .CP(clk), .CD(n18256), .Q(Poly15[55])
         );
  CFD2QXL \Poly14_reg[285]  ( .D(n10120), .CP(clk), .CD(n18310), .Q(
        Poly14[285]) );
  CFD2QXL \Poly13_reg[527]  ( .D(n10533), .CP(clk), .CD(n18274), .Q(
        Poly13[527]) );
  CFD2QXL \Poly13_reg[520]  ( .D(n10540), .CP(clk), .CD(n18287), .Q(
        Poly13[520]) );
  CFD2QXL \Poly11_reg[85]  ( .D(n11104), .CP(clk), .CD(n18257), .Q(Poly11[85])
         );
  CFD2QXL \Poly11_reg[78]  ( .D(n11111), .CP(clk), .CD(n18257), .Q(Poly11[78])
         );
  CFD2QXL \Poly5_reg[114]  ( .D(n11412), .CP(clk), .CD(n18258), .Q(Poly5[114])
         );
  CFD2QXL \Poly15_reg[57]  ( .D(n9580), .CP(clk), .CD(n18345), .Q(Poly15[57])
         );
  CFD2QXL \Poly2_reg[64]  ( .D(n8946), .CP(clk), .CD(n18378), .Q(Poly2[64]) );
  CFD2QXL \Poly2_reg[68]  ( .D(n8942), .CP(clk), .CD(n18379), .Q(Poly2[68]) );
  CFD2QXL \Poly12_reg[126]  ( .D(n10406), .CP(clk), .CD(n18294), .Q(
        Poly12[126]) );
  CFD2QXL \Poly11_reg[80]  ( .D(n11109), .CP(clk), .CD(n18257), .Q(Poly11[80])
         );
  CFD2QXL \Poly12_reg[117]  ( .D(n10415), .CP(clk), .CD(n18295), .Q(
        Poly12[117]) );
  CFD2QXL \Poly12_reg[114]  ( .D(n10418), .CP(clk), .CD(n18292), .Q(
        Poly12[114]) );
  CFD2QXL \Poly10_reg[38]  ( .D(n11065), .CP(clk), .CD(n18400), .Q(Poly10[38])
         );
  CFD2QXL \Poly12_reg[125]  ( .D(n10407), .CP(clk), .CD(n18297), .Q(
        Poly12[125]) );
  CFD2QXL \Poly11_reg[81]  ( .D(n11108), .CP(clk), .CD(n18257), .Q(Poly11[81])
         );
  CFD2QXL \Poly0_reg[143]  ( .D(n9434), .CP(clk), .CD(n18356), .Q(
        poly0_shifted[161]) );
  CFD2QXL \Poly0_reg[161]  ( .D(n9416), .CP(clk), .CD(n18356), .Q(Poly0[161])
         );
  CFD2QXL \Poly2_reg[59]  ( .D(n8951), .CP(clk), .CD(n18380), .Q(Poly2[59]) );
  CFD2QXL \Poly11_reg[76]  ( .D(n11113), .CP(clk), .CD(n18257), .Q(Poly11[76])
         );
  CFD2QXL \Poly4_reg[48]  ( .D(n8808), .CP(clk), .CD(n18389), .Q(Poly4[48]) );
  CFD2QXL \Poly4_reg[44]  ( .D(n8812), .CP(clk), .CD(n18386), .Q(Poly4[44]) );
  CFD2QXL \Poly4_reg[45]  ( .D(n8811), .CP(clk), .CD(n18389), .Q(Poly4[45]) );
  CFD2QXL \dataselector_reg[5]  ( .D(n8790), .CP(clk), .CD(n18388), .Q(
        dataselector[5]) );
  CFD2QXL \Poly11_reg[74]  ( .D(n11115), .CP(clk), .CD(n18262), .Q(Poly11[74])
         );
  CFD2QXL \Poly4_reg[46]  ( .D(n8810), .CP(clk), .CD(n18389), .Q(Poly4[46]) );
  CFD2QXL \Poly4_reg[49]  ( .D(n8807), .CP(clk), .CD(n18389), .Q(Poly4[49]) );
  CFD2QXL \dataselector_reg[8]  ( .D(n8787), .CP(clk), .CD(n18387), .Q(
        dataselector[8]) );
  CFD2QXL \Poly2_reg[66]  ( .D(n8944), .CP(clk), .CD(n18378), .Q(Poly2[66]) );
  CFD2QX1 \scrambler_reg[25]  ( .D(n8725), .CP(clk), .CD(n18401), .Q(
        scrambler[25]) );
  CFD2QXL \Poly4_reg[47]  ( .D(n8809), .CP(clk), .CD(n18389), .Q(Poly4[47]) );
  CFD2QXL \Poly2_reg[67]  ( .D(n8943), .CP(clk), .CD(n18378), .Q(Poly2[67]) );
  CFD2QX1 \dataselector_reg[61]  ( .D(n8734), .CP(clk), .CD(n18386), .Q(
        dataselector[61]) );
  CFD2QXL \dataselector_reg[31]  ( .D(n8764), .CP(clk), .CD(n18388), .Q(
        dataselector[31]) );
  CFD2QX1 \Poly4_reg[58]  ( .D(n8798), .CP(clk), .CD(n18385), .Q(Poly4[58]) );
  CFD2QXL \Poly6_reg[52]  ( .D(n9641), .CP(clk), .CD(n18343), .Q(Poly6[52]) );
  CFD2QX1 \dataselector_reg[57]  ( .D(n8738), .CP(clk), .CD(n18386), .Q(
        dataselector[57]) );
  CFD2QXL \Poly11_reg[79]  ( .D(n11110), .CP(clk), .CD(n18257), .Q(Poly11[79])
         );
  CFD2QXL \Poly11_reg[82]  ( .D(n11107), .CP(clk), .CD(n18257), .Q(Poly11[82])
         );
  CFD2QXL \dataselector_reg[47]  ( .D(n8748), .CP(clk), .CD(n18402), .Q(
        dataselector[47]) );
  CFD2QXL \dataselector_reg[53]  ( .D(n8742), .CP(clk), .CD(n18387), .Q(
        dataselector[53]) );
  CFD2QX1 \dataselector_reg[60]  ( .D(n8735), .CP(clk), .CD(n18402), .Q(
        dataselector[60]) );
  CFD2QXL \scrambler_reg[27]  ( .D(n8727), .CP(clk), .CD(n18401), .Q(
        scrambler[27]) );
  CFD2QXL \scrambler_reg[16]  ( .D(n8716), .CP(clk), .CD(n18257), .Q(
        scrambler[16]) );
  CFD2QX1 \dataselector_reg[25]  ( .D(n8770), .CP(clk), .CD(n18402), .Q(
        dataselector[25]) );
  CFD2QXL \Poly11_reg[83]  ( .D(n11106), .CP(clk), .CD(n18257), .Q(Poly11[83])
         );
  CFD2QXL \Poly2_reg[65]  ( .D(n8945), .CP(clk), .CD(n18392), .Q(Poly2[65]) );
  CFD2QXL \Poly11_reg[84]  ( .D(n11105), .CP(clk), .CD(n18257), .Q(Poly11[84])
         );
  CFD2QXL \scrambler_reg[30]  ( .D(n8730), .CP(clk), .CD(n18401), .Q(
        scrambler[30]) );
  CFD2QXL \scrambler_reg[19]  ( .D(n8719), .CP(clk), .CD(n18257), .Q(
        scrambler[19]) );
  CFD2QXL \scrambler_reg[31]  ( .D(n8731), .CP(clk), .CD(n18257), .Q(
        scrambler[31]) );
  CFD2QXL \scrambler_reg[29]  ( .D(n8729), .CP(clk), .CD(n18257), .Q(
        scrambler[29]) );
  CFD2QXL \Poly4_reg[55]  ( .D(n8801), .CP(clk), .CD(n18256), .Q(Poly4[55]) );
  CFD2QX2 \scrambler_reg[20]  ( .D(n8720), .CP(clk), .CD(n18257), .Q(
        scrambler[20]) );
  CFD2QX1 \Poly4_reg[51]  ( .D(n8805), .CP(clk), .CD(n18389), .Q(Poly4[51]) );
  CFD2QXL \dataselector_reg[1]  ( .D(n8794), .CP(clk), .CD(n18389), .Q(
        dataselector[1]) );
  CFD2QXL \polydata_reg[0]  ( .D(n8684), .CP(clk), .CD(n18257), .Q(polydata[0]) );
  CFD2QXL \polydata_reg[5]  ( .D(n8689), .CP(clk), .CD(n18257), .Q(polydata[5]) );
  CFD2QXL \polydata_reg[4]  ( .D(n8688), .CP(clk), .CD(n18401), .Q(polydata[4]) );
  CFD2QX1 \Poly4_reg[53]  ( .D(n8803), .CP(clk), .CD(n18385), .Q(Poly4[53]) );
  CFD2QXL \scrambler_reg[23]  ( .D(n8723), .CP(clk), .CD(n18401), .Q(
        scrambler[23]) );
  CIVDX1 U8718 ( .A(n15306), .Z0(n14935), .Z1(n17770) );
  CNR2X1 U8719 ( .A(n15349), .B(n13958), .Z(n15043) );
  CAN2X1 U8720 ( .A(n13878), .B(n15583), .Z(n18046) );
  CNR2X1 U8721 ( .A(n12059), .B(n12058), .Z(n12060) );
  CNR2X2 U8722 ( .A(n12596), .B(dataselector[5]), .Z(n12073) );
  CANR1XL U8723 ( .A(entrophy[27]), .B(n15052), .C(n14641), .Z(n14642) );
  COND1XL U8724 ( .A(n15044), .B(n14640), .C(n14866), .Z(n14641) );
  CND2X1 U8725 ( .A(n12092), .B(n13780), .Z(n12108) );
  CND2X1 U8726 ( .A(n13781), .B(n18244), .Z(n12074) );
  CND3X2 U8727 ( .A(n12091), .B(n12385), .C(n12596), .Z(n12104) );
  CIVX2 U8728 ( .A(n14887), .Z(n12534) );
  CANR1X1 U8729 ( .A(entrophy[19]), .B(n17812), .C(n14861), .Z(n14862) );
  CNR2X1 U8730 ( .A(n14633), .B(n14632), .Z(n14669) );
  CND3XL U8731 ( .A(n15160), .B(n14085), .C(n12214), .Z(n14218) );
  CNR3X1 U8732 ( .A(n13953), .B(n13952), .C(n13951), .Z(n13954) );
  CND3XL U8733 ( .A(n15143), .B(n13949), .C(n13948), .Z(n13953) );
  CNR2X1 U8734 ( .A(n14472), .B(n14908), .Z(n14823) );
  CND2IX1 U8735 ( .B(n12278), .A(n12209), .Z(n12649) );
  CNIVX2 U8736 ( .A(n15319), .Z(n11974) );
  CNR3XL U8737 ( .A(n14538), .B(n17763), .C(n14561), .Z(n14539) );
  CNIVX4 U8738 ( .A(n12111), .Z(n16864) );
  CND2X1 U8739 ( .A(n15256), .B(entrophy[23]), .Z(n14846) );
  CNR2X1 U8740 ( .A(n12534), .B(n14395), .Z(n15249) );
  CAN2X1 U8741 ( .A(n15206), .B(n12216), .Z(n17787) );
  CANR1XL U8742 ( .A(n17805), .B(n14966), .C(n11969), .Z(n12444) );
  CIVX2 U8743 ( .A(n12241), .Z(n12092) );
  CND2X1 U8744 ( .A(addr[1]), .B(n12166), .Z(n12404) );
  CND2X1 U8745 ( .A(addr[1]), .B(addr[0]), .Z(n12243) );
  CND2X1 U8746 ( .A(addr[6]), .B(n12151), .Z(n12191) );
  CND2IX1 U8747 ( .B(n12243), .A(n12209), .Z(n12680) );
  CND2IX1 U8748 ( .B(n12200), .A(addr[6]), .Z(n12269) );
  CNR2IX1 U8749 ( .B(n15302), .A(n14797), .Z(n15119) );
  CND2IX1 U8750 ( .B(n12165), .A(dataselector[53]), .Z(n12241) );
  CANR1X1 U8751 ( .A(n12216), .B(n14144), .C(n14143), .Z(n14145) );
  COND1XL U8752 ( .A(n14991), .B(n14990), .C(n15145), .Z(n14992) );
  CND2IX1 U8753 ( .B(n12173), .A(n14393), .Z(n14796) );
  CIVX2 U8754 ( .A(n12598), .Z(n13511) );
  CNIVX4 U8755 ( .A(n13137), .Z(n17603) );
  CIVX2 U8756 ( .A(n15648), .Z(n17640) );
  CNIVX4 U8757 ( .A(n12361), .Z(n17977) );
  CNR2X2 U8758 ( .A(n12649), .B(n12648), .Z(n18209) );
  CNR2X2 U8759 ( .A(n18209), .B(n16947), .Z(n17359) );
  CNIVX2 U8760 ( .A(n12279), .Z(n14441) );
  CIVDX1 U8761 ( .A(n12382), .Z0(n13443), .Z1(n13840) );
  CNIVX4 U8762 ( .A(n13146), .Z(n17955) );
  CIVX2 U8763 ( .A(n17076), .Z(n18048) );
  CNIVX4 U8764 ( .A(n12611), .Z(n17595) );
  CNIVX4 U8765 ( .A(n12270), .Z(n17990) );
  CNIVX3 U8766 ( .A(n17564), .Z(n18018) );
  CNR2IX1 U8767 ( .B(Poly12[119]), .A(n17495), .Z(n17994) );
  COND1X1 U8768 ( .A(n17774), .B(n15330), .C(datain[1]), .Z(n14933) );
  CNIVX1 U8769 ( .A(n17805), .Z(n11972) );
  CIVX4 U8770 ( .A(n12266), .Z(n17714) );
  CIVX2 U8771 ( .A(n16248), .Z(n18206) );
  CNIVX4 U8772 ( .A(n12212), .Z(n18044) );
  CAN2X1 U8773 ( .A(n17826), .B(lfsrdin[29]), .Z(n18228) );
  CAN2X1 U8774 ( .A(n12396), .B(n13266), .Z(n13782) );
  CENX1 U8775 ( .A(dataselector[63]), .B(n18253), .Z(n18239) );
  CIVX8 U8776 ( .A(n17826), .Z(n18234) );
  CNR2X2 U8777 ( .A(n17317), .B(n15960), .Z(n15671) );
  CNIVX4 U8778 ( .A(n13879), .Z(n17525) );
  CIVX4 U8779 ( .A(n18099), .Z(n17741) );
  CNIVX4 U8780 ( .A(n12995), .Z(n18002) );
  CNIVX4 U8781 ( .A(n13239), .Z(n17969) );
  CIVX2 U8782 ( .A(n12381), .Z(n17062) );
  CND2X2 U8783 ( .A(n12763), .B(n13227), .Z(n15880) );
  CIVX4 U8784 ( .A(n15648), .Z(n17620) );
  CAN2X1 U8785 ( .A(n17829), .B(lfsrdin[19]), .Z(n18176) );
  CIVX8 U8786 ( .A(n15648), .Z(n17755) );
  CIVDX1 U8787 ( .A(n12914), .Z0(n12915), .Z1(n14166) );
  CIVX4 U8788 ( .A(n13663), .Z(n17750) );
  CIVX2 U8789 ( .A(n15648), .Z(n17560) );
  CNIVX2 U8790 ( .A(n12273), .Z(n12006) );
  CIVDX2 U8791 ( .A(n12296), .Z0(n11999), .Z1(n12000) );
  CND2X1 U8792 ( .A(n17200), .B(n17826), .Z(n18196) );
  CIVX2 U8793 ( .A(n14944), .Z(n17832) );
  CND3XL U8794 ( .A(n14370), .B(n14217), .C(n14888), .Z(n14706) );
  CIVX2 U8795 ( .A(n16139), .Z(n18248) );
  CIVX2 U8796 ( .A(n12553), .Z(n14788) );
  CAN2X2 U8797 ( .A(n17495), .B(lfsrdin[18]), .Z(n18210) );
  CAN2X1 U8798 ( .A(n17495), .B(lfsrdin[27]), .Z(n18099) );
  CND2X2 U8799 ( .A(dataselector[31]), .B(n12085), .Z(n12102) );
  CIVX4 U8800 ( .A(n12106), .Z(n12114) );
  CND2IX1 U8801 ( .B(addr[1]), .A(n12166), .Z(n12278) );
  CND2X1 U8802 ( .A(addr[3]), .B(n12159), .Z(n12277) );
  CNR2X2 U8803 ( .A(n12953), .B(n18184), .Z(n14159) );
  CND2X2 U8804 ( .A(n12680), .B(n17959), .Z(n13227) );
  CIVX8 U8805 ( .A(n11975), .Z(n13878) );
  COAN1X1 U8806 ( .A(n12261), .B(n12269), .C(n17495), .Z(n11975) );
  CNR3XL U8807 ( .A(n14452), .B(n14644), .C(n14977), .Z(n14481) );
  CND3X1 U8808 ( .A(n12545), .B(n12544), .C(n12543), .Z(n8708) );
  CND2IX1 U8809 ( .B(n12529), .A(n12528), .Z(n12545) );
  COND1XL U8810 ( .A(n16565), .B(n16745), .C(n16744), .Z(n9601) );
  CNIVX1 U8811 ( .A(n18257), .Z(n18254) );
  CNIVX1 U8812 ( .A(n18257), .Z(n18255) );
  CND4X1 U8813 ( .A(n12063), .B(n12062), .C(n12061), .D(n12060), .Z(n8722) );
  CNIVX1 U8814 ( .A(n18257), .Z(n18256) );
  CNR2X1 U8815 ( .A(n12110), .B(n12112), .Z(n12086) );
  CNR2X1 U8816 ( .A(n12110), .B(n12114), .Z(n12111) );
  CIVX1 U8817 ( .A(n15335), .Z(n11527) );
  CANR2X1 U8818 ( .A(n15046), .B(n15354), .C(n15045), .D(n11527), .Z(n15051)
         );
  CND2IX1 U8819 ( .B(n15059), .A(n15060), .Z(n15067) );
  CANR3X1 U8820 ( .A(n15348), .B(datain[1]), .C(n14233), .D(n14232), .Z(n11528) );
  CAN4X1 U8821 ( .A(n15071), .B(n15172), .C(n15096), .D(n15142), .Z(n11529) );
  COND4CX1 U8822 ( .A(n11528), .B(n11529), .C(n15334), .D(n15170), .Z(n14234)
         );
  COND1XL U8823 ( .A(n15299), .B(n14966), .C(n14890), .Z(n11530) );
  CNR2X1 U8824 ( .A(n15091), .B(n11530), .Z(n11531) );
  CND3XL U8825 ( .A(n14590), .B(n13949), .C(n11531), .Z(n12441) );
  CND2IX1 U8826 ( .B(Poly2[65]), .A(n16947), .Z(n13754) );
  CIVX2 U8827 ( .A(n18039), .Z(n12007) );
  CND2X1 U8828 ( .A(poly5_shifted[36]), .B(n17640), .Z(n11532) );
  CMXI2X1 U8829 ( .A0(poly5_shifted[50]), .A1(n12004), .S(n12942), .Z(n11533)
         );
  CND2X1 U8830 ( .A(n11532), .B(n11533), .Z(n11490) );
  CND2X1 U8831 ( .A(poly5_shifted[86]), .B(n17215), .Z(n11534) );
  CMXI2X1 U8832 ( .A0(Poly5[86]), .A1(n18034), .S(n17045), .Z(n11535) );
  CND2X1 U8833 ( .A(n11534), .B(n11535), .Z(n11440) );
  CIVX1 U8834 ( .A(n14982), .Z(n11536) );
  CAN3X1 U8835 ( .A(n14416), .B(n14683), .C(n11536), .Z(n13948) );
  CND2X1 U8836 ( .A(entrophy[11]), .B(n14826), .Z(n11537) );
  CND3XL U8837 ( .A(n11537), .B(n14684), .C(n14845), .Z(n12223) );
  COND3X1 U8838 ( .A(n14967), .B(n14644), .C(n14643), .D(n14642), .Z(n14658)
         );
  CANR4CX1 U8839 ( .A(n14838), .B(n14129), .C(n15220), .D(n13959), .Z(n11538)
         );
  COND3X1 U8840 ( .A(n14788), .B(n14705), .C(n13960), .D(n11538), .Z(n13966)
         );
  CND2IX1 U8841 ( .B(Poly6[54]), .A(n17317), .Z(n16959) );
  CIVX1 U8842 ( .A(n14690), .Z(n11539) );
  CNR2X1 U8843 ( .A(n14473), .B(n14807), .Z(n11540) );
  CNR8X1 U8844 ( .A(n11539), .B(n12521), .C(n14093), .D(n12536), .E(n15017), 
        .F(n15205), .G(n11540), .H(n15144), .Z(n12529) );
  CANR2X1 U8845 ( .A(poly1_shifted[259]), .B(n16872), .C(poly2_shifted[25]), 
        .D(n16843), .Z(n11541) );
  CANR2X1 U8846 ( .A(n16864), .B(poly0_shifted[163]), .C(n16729), .D(n16852), 
        .Z(n11542) );
  CAN4X1 U8847 ( .A(n11541), .B(n11542), .C(n16730), .D(n16731), .Z(n16737) );
  COND1XL U8848 ( .A(poly0_shifted[219]), .B(n18099), .C(n18098), .Z(n11543)
         );
  CND2X1 U8849 ( .A(n18119), .B(Poly0[219]), .Z(n11544) );
  COND1XL U8850 ( .A(n18119), .B(n11543), .C(n11544), .Z(n9358) );
  COND1XL U8851 ( .A(Poly5[123]), .B(Poly5[101]), .C(n17634), .Z(n11545) );
  CMXI2X1 U8852 ( .A0(Poly5[115]), .A1(n18176), .S(n15574), .Z(n11546) );
  COND4CX1 U8853 ( .A(Poly5[101]), .B(Poly5[123]), .C(n11545), .D(n11546), .Z(
        n11411) );
  CENX1 U8854 ( .A(Poly8[88]), .B(Poly8[73]), .Z(n11547) );
  CMXI2X1 U8855 ( .A0(n11999), .A1(Poly8[87]), .S(n17750), .Z(n11548) );
  COND1XL U8856 ( .A(n17160), .B(n11547), .C(n11548), .Z(n11314) );
  COND1XL U8857 ( .A(poly10_shifted[40]), .B(n18142), .C(n18141), .Z(n11549)
         );
  CND2X1 U8858 ( .A(n17411), .B(Poly10[40]), .Z(n11550) );
  COND1XL U8859 ( .A(n17411), .B(n11549), .C(n11550), .Z(n11063) );
  CNR2X1 U8860 ( .A(n16753), .B(Poly2[42]), .Z(n11551) );
  CNR2X1 U8861 ( .A(n18034), .B(n11551), .Z(n11552) );
  CANR2X1 U8862 ( .A(n17306), .B(Poly2[54]), .C(Poly2[42]), .D(n13553), .Z(
        n11553) );
  COND1XL U8863 ( .A(n17306), .B(n11552), .C(n11553), .Z(n8956) );
  CND2X1 U8864 ( .A(poly5_shifted[35]), .B(n17238), .Z(n11554) );
  CMXI2X1 U8865 ( .A0(poly5_shifted[49]), .A1(n18053), .S(n12942), .Z(n11555)
         );
  CND2X1 U8866 ( .A(n11554), .B(n11555), .Z(n11491) );
  CAOR2X1 U8867 ( .A(n17495), .B(scrambler[3]), .C(n14976), .D(n15045), .Z(
        n12486) );
  CNR2IX1 U8868 ( .B(n17767), .A(n14960), .Z(n15312) );
  CNR2X1 U8869 ( .A(n14982), .B(n14091), .Z(n11556) );
  COND11X1 U8870 ( .A(n14395), .B(n14968), .C(n14887), .D(n11556), .Z(n14092)
         );
  CND4X1 U8871 ( .A(n15329), .B(n15097), .C(n12222), .D(n15252), .Z(n11557) );
  CNR3X1 U8872 ( .A(n12223), .B(n15286), .C(n11557), .Z(n12230) );
  CND3XL U8873 ( .A(n12038), .B(n12037), .C(n17763), .Z(n12039) );
  CNR2X2 U8874 ( .A(n14963), .B(n15218), .Z(n11971) );
  CIVX2 U8875 ( .A(n11971), .Z(n11970) );
  CANR2X1 U8876 ( .A(n16863), .B(Poly8[68]), .C(n16850), .D(Poly5[122]), .Z(
        n11558) );
  CANR2X1 U8877 ( .A(Poly3[57]), .B(n16844), .C(n16750), .D(n16840), .Z(n11559) );
  CAN4X1 U8878 ( .A(n11558), .B(n11559), .C(n16751), .D(n16752), .Z(n16765) );
  COND1XL U8879 ( .A(n17163), .B(n14944), .C(n12596), .Z(n11560) );
  CANR1XL U8880 ( .A(dataselector[8]), .B(n16410), .C(n11560), .Z(n11561) );
  COND1XL U8881 ( .A(n17830), .B(dataselector[61]), .C(n17535), .Z(n11562) );
  CANR1XL U8882 ( .A(n17830), .B(dataselector[61]), .C(n11562), .Z(n11563) );
  CMXI2X1 U8883 ( .A0(n11561), .A1(dataselector[1]), .S(n11563), .Z(n8787) );
  CIVX1 U8884 ( .A(n15673), .Z(n11564) );
  CIVX1 U8885 ( .A(n15672), .Z(n11565) );
  CANR2X1 U8886 ( .A(poly0_shifted[161]), .B(n11564), .C(Poly0[161]), .D(
        n11565), .Z(n11566) );
  COND1XL U8887 ( .A(n17316), .B(n17711), .C(n11566), .Z(n9416) );
  CND2X1 U8888 ( .A(poly5_shifted[123]), .B(n17998), .Z(n11567) );
  CMXI2X1 U8889 ( .A0(Poly5[123]), .A1(n18099), .S(n17031), .Z(n11568) );
  CND2X1 U8890 ( .A(n11567), .B(n11568), .Z(n11403) );
  CEOX1 U8891 ( .A(Poly2[64]), .B(Poly2[57]), .Z(n11569) );
  CND2X1 U8892 ( .A(n11569), .B(n13553), .Z(n11570) );
  COND1XL U8893 ( .A(n16753), .B(n11569), .C(n11987), .Z(n11571) );
  CMXI2X1 U8894 ( .A0(n11571), .A1(Poly2[69]), .S(n17696), .Z(n11572) );
  CND2X1 U8895 ( .A(n11570), .B(n11572), .Z(n8941) );
  COND1XL U8896 ( .A(poly0_shifted[205]), .B(n18219), .C(n18156), .Z(n11573)
         );
  CND2X1 U8897 ( .A(n18119), .B(Poly0[205]), .Z(n11574) );
  COND1XL U8898 ( .A(n18119), .B(n11573), .C(n11574), .Z(n9372) );
  CND2X1 U8899 ( .A(n18050), .B(Poly15[16]), .Z(n11575) );
  CND3XL U8900 ( .A(n17317), .B(n14322), .C(n11575), .Z(n11576) );
  CNR2X1 U8901 ( .A(n11575), .B(n14323), .Z(n11577) );
  CANR1XL U8902 ( .A(Poly15[31]), .B(n18044), .C(n11577), .Z(n11578) );
  COND4CX1 U8903 ( .A(n17188), .B(n11576), .C(n18044), .D(n11578), .Z(n9606)
         );
  COND1XL U8904 ( .A(poly0_shifted[93]), .B(n18228), .C(n18227), .Z(n11579) );
  CND2X1 U8905 ( .A(n12291), .B(poly0_shifted[111]), .Z(n11580) );
  COND1XL U8906 ( .A(n12291), .B(n11579), .C(n11580), .Z(n9484) );
  COND1XL U8907 ( .A(poly5_shifted[22]), .B(n18034), .C(n18088), .Z(n11581) );
  CND2X1 U8908 ( .A(n17932), .B(poly5_shifted[36]), .Z(n11582) );
  COND1XL U8909 ( .A(n17932), .B(n11581), .C(n11582), .Z(n11504) );
  CND2X1 U8910 ( .A(poly5_shifted[43]), .B(n17238), .Z(n11583) );
  CMXI2X1 U8911 ( .A0(poly5_shifted[57]), .A1(n16381), .S(n12942), .Z(n11584)
         );
  CND2X1 U8912 ( .A(n11583), .B(n11584), .Z(n11483) );
  CANR1XL U8913 ( .A(Poly10[0]), .B(Poly10[38]), .C(n17160), .Z(n11585) );
  CANR4CX1 U8914 ( .A(Poly10[0]), .B(Poly10[38]), .C(n11585), .D(n13028), .Z(
        n11586) );
  CMXI2X1 U8915 ( .A0(n13759), .A1(n11586), .S(n13782), .Z(n11091) );
  CANR1XL U8916 ( .A(n15206), .B(datain[2]), .C(n15311), .Z(n14892) );
  CND2IX1 U8917 ( .B(n15219), .A(n14669), .Z(n14650) );
  CIVX1 U8918 ( .A(n15216), .Z(n11587) );
  CND4X1 U8919 ( .A(n15217), .B(n15214), .C(n15215), .D(n11587), .Z(n15222) );
  CND2IX1 U8920 ( .B(n15168), .A(n15169), .Z(n11588) );
  CAN4X1 U8921 ( .A(n15165), .B(n15167), .C(n15166), .D(n11588), .Z(n15174) );
  CNR2X1 U8922 ( .A(n11972), .B(n14886), .Z(n11589) );
  CND2X1 U8923 ( .A(n14887), .B(n11589), .Z(n11590) );
  CND4X1 U8924 ( .A(n15287), .B(n14888), .C(n15115), .D(n11590), .Z(n14889) );
  CIVX1 U8925 ( .A(n14977), .Z(n11591) );
  CND4X1 U8926 ( .A(n14638), .B(n14639), .C(n15097), .D(n15142), .Z(n11592) );
  CND3XL U8927 ( .A(n14658), .B(n11591), .C(n11592), .Z(n14677) );
  CND2IX1 U8928 ( .B(Poly15[46]), .A(n17755), .Z(n13940) );
  CNR3XL U8929 ( .A(n14936), .B(n15112), .C(n14966), .Z(n11593) );
  COND1XL U8930 ( .A(n14558), .B(n17763), .C(n14557), .Z(n11594) );
  CANR3X1 U8931 ( .A(n17812), .B(entrophy[5]), .C(n11593), .D(n11594), .Z(
        n14564) );
  CANR2X1 U8932 ( .A(poly12_shifted[88]), .B(n16853), .C(poly13_shifted[25]), 
        .D(n16875), .Z(n11595) );
  CANR2X1 U8933 ( .A(Poly15[47]), .B(n12067), .C(poly12_shifted[122]), .D(
        n16855), .Z(n11596) );
  CAN4X1 U8934 ( .A(n11595), .B(n11596), .C(n16830), .D(n16831), .Z(n16832) );
  CIVX1 U8935 ( .A(n15309), .Z(n11597) );
  COND11X1 U8936 ( .A(n12460), .B(n12501), .C(n12461), .D(n15220), .Z(n11598)
         );
  COND1XL U8937 ( .A(n14947), .B(n11597), .C(n11598), .Z(n12462) );
  CENX1 U8938 ( .A(n16385), .B(Poly7[409]), .Z(n11599) );
  CNR2X1 U8939 ( .A(n11599), .B(n17959), .Z(n11600) );
  CANR1XL U8940 ( .A(n16410), .B(dataselector[5]), .C(n11600), .Z(n11601) );
  COND1XL U8941 ( .A(n11991), .B(n14944), .C(n11601), .Z(n8790) );
  COND1XL U8942 ( .A(poly14_shifted[289]), .B(n12020), .C(n18123), .Z(n11602)
         );
  CND2X1 U8943 ( .A(n17444), .B(Poly14[289]), .Z(n11603) );
  COND1XL U8944 ( .A(n17444), .B(n11602), .C(n11603), .Z(n10116) );
  COND1XL U8945 ( .A(poly0_shifted[218]), .B(n18095), .C(n18094), .Z(n11604)
         );
  CND2X1 U8946 ( .A(n18119), .B(Poly0[218]), .Z(n11605) );
  COND1XL U8947 ( .A(n18119), .B(n11604), .C(n11605), .Z(n9359) );
  COND1XL U8948 ( .A(poly0_shifted[214]), .B(n14487), .C(n18088), .Z(n11606)
         );
  CND2X1 U8949 ( .A(n18119), .B(Poly0[214]), .Z(n11607) );
  COND1XL U8950 ( .A(n18119), .B(n11606), .C(n11607), .Z(n9363) );
  COND1XL U8951 ( .A(poly0_shifted[213]), .B(n18241), .C(n18085), .Z(n11608)
         );
  CND2X1 U8952 ( .A(n18119), .B(Poly0[213]), .Z(n11609) );
  COND1XL U8953 ( .A(n18119), .B(n11608), .C(n11609), .Z(n9364) );
  COND1XL U8954 ( .A(n13522), .B(poly0_shifted[209]), .C(n18193), .Z(n11610)
         );
  CND2X1 U8955 ( .A(n18119), .B(Poly0[209]), .Z(n11611) );
  COND1XL U8956 ( .A(n18119), .B(n11610), .C(n11611), .Z(n9368) );
  COND1XL U8957 ( .A(poly0_shifted[216]), .B(n13994), .C(n18091), .Z(n11612)
         );
  CND2X1 U8958 ( .A(n18119), .B(Poly0[216]), .Z(n11613) );
  COND1XL U8959 ( .A(n18119), .B(n11612), .C(n11613), .Z(n9361) );
  COND1XL U8960 ( .A(poly10_shifted[39]), .B(n18138), .C(n18137), .Z(n11614)
         );
  CND2X1 U8961 ( .A(n17411), .B(Poly10[39]), .Z(n11615) );
  COND1XL U8962 ( .A(n17411), .B(n11614), .C(n11615), .Z(n11064) );
  COND1XL U8963 ( .A(poly2_shifted[25]), .B(n17934), .C(n18196), .Z(n11616) );
  CND2X1 U8964 ( .A(n12211), .B(Poly2[25]), .Z(n11617) );
  COND1XL U8965 ( .A(n12211), .B(n11616), .C(n11617), .Z(n8985) );
  CMXI2X1 U8966 ( .A0(n17994), .A1(poly12_shifted[24]), .S(n12997), .Z(n11618)
         );
  COND1XL U8967 ( .A(n12997), .B(n17163), .C(n11618), .Z(n10524) );
  CND3XL U8968 ( .A(Poly11[21]), .B(n17628), .C(n17317), .Z(n11619) );
  CNR2X1 U8969 ( .A(Poly11[21]), .B(n15246), .Z(n11620) );
  CANR1XL U8970 ( .A(n17683), .B(Poly11[36]), .C(n11620), .Z(n11621) );
  COND4CX1 U8971 ( .A(n12005), .B(n11619), .C(n17683), .D(n11621), .Z(n11153)
         );
  CMX2GX1 U8972 ( .GN(n18099), .A0(n13453), .A1(n13452), .S(Poly6[17]), .Z(
        n11622) );
  CND2X1 U8973 ( .A(n13840), .B(Poly6[27]), .Z(n11623) );
  COND1XL U8974 ( .A(n11622), .B(n13840), .C(n11623), .Z(n9666) );
  COND1XL U8975 ( .A(poly13_shifted[493]), .B(n18219), .C(n18156), .Z(n11624)
         );
  CND2X1 U8976 ( .A(n17491), .B(poly13_shifted[507]), .Z(n11625) );
  COND1XL U8977 ( .A(n17491), .B(n11624), .C(n11625), .Z(n10567) );
  COND1XL U8978 ( .A(poly9_shifted[60]), .B(n12007), .C(n18224), .Z(n11626) );
  CND2X1 U8979 ( .A(n13351), .B(poly9_shifted[71]), .Z(n11627) );
  COND1XL U8980 ( .A(n13351), .B(n11626), .C(n11627), .Z(n11245) );
  CIVX1 U8981 ( .A(n15571), .Z(n11628) );
  COND1XL U8982 ( .A(n14754), .B(n11628), .C(n18117), .Z(n11629) );
  CND2X1 U8983 ( .A(n15378), .B(poly5_shifted[52]), .Z(n11630) );
  COND1XL U8984 ( .A(n15378), .B(n11629), .C(n11630), .Z(n11488) );
  COND1XL U8985 ( .A(poly3_shifted[42]), .B(n12013), .C(n18147), .Z(n11631) );
  CND2X1 U8986 ( .A(n17262), .B(Poly3[42]), .Z(n11632) );
  COND1XL U8987 ( .A(n17262), .B(n11631), .C(n11632), .Z(n8898) );
  CMXI2X1 U8988 ( .A0(Poly5[93]), .A1(n18228), .S(n17045), .Z(n11633) );
  COND1XL U8989 ( .A(Poly5[114]), .B(Poly5[79]), .C(n17705), .Z(n11634) );
  COND4CX1 U8990 ( .A(Poly5[79]), .B(Poly5[114]), .C(n11634), .D(n11633), .Z(
        n11433) );
  CANR2X1 U8991 ( .A(n12299), .B(poly1_shifted[60]), .C(poly1_shifted[49]), 
        .D(n16947), .Z(n11635) );
  COND1XL U8992 ( .A(n12299), .B(n17173), .C(n11635), .Z(n9308) );
  CND2X1 U8993 ( .A(poly5_shifted[37]), .B(n18234), .Z(n11636) );
  CMXI2X1 U8994 ( .A0(poly5_shifted[51]), .A1(n11988), .S(n12942), .Z(n11637)
         );
  CND2X1 U8995 ( .A(n11636), .B(n11637), .Z(n11489) );
  CMX2GX1 U8996 ( .GN(n18034), .A0(n13468), .A1(n13467), .S(Poly6[12]), .Z(
        n11638) );
  CND2X1 U8997 ( .A(n14310), .B(Poly6[22]), .Z(n11639) );
  COND1XL U8998 ( .A(n11638), .B(n14310), .C(n11639), .Z(n9671) );
  COND3X1 U8999 ( .A(n15256), .B(entrophy[4]), .C(n12444), .D(n14369), .Z(
        n12472) );
  CND3XL U9000 ( .A(n14797), .B(entrophy[26]), .C(n14392), .Z(n11640) );
  CND3XL U9001 ( .A(n11640), .B(n12053), .C(n12052), .Z(n11641) );
  CND2X1 U9002 ( .A(n11641), .B(n15220), .Z(n12056) );
  CND8X1 U9003 ( .A(n14704), .B(n15140), .C(n14986), .D(n15070), .E(n14227), 
        .F(n14228), .G(n14229), .H(n14689), .Z(n11642) );
  CND2X1 U9004 ( .A(n14234), .B(n11642), .Z(n14235) );
  COND1XL U9005 ( .A(n12018), .B(n14453), .C(n14893), .Z(n14418) );
  CNR2IX1 U9006 ( .B(n13493), .A(Poly6[52]), .Z(n13815) );
  CND2IX1 U9007 ( .B(n12256), .A(n17538), .Z(n17310) );
  CANR2X1 U9008 ( .A(poly8_shifted[50]), .B(n16864), .C(Poly8[73]), .D(n16855), 
        .Z(n11643) );
  CANR2X1 U9009 ( .A(n16854), .B(poly1_shifted[315]), .C(poly8_shifted[77]), 
        .D(n16866), .Z(n11644) );
  CAN4X1 U9010 ( .A(n11643), .B(n11644), .C(n16806), .D(n16807), .Z(n16813) );
  CANR1XL U9011 ( .A(entrophy[2]), .B(n15330), .C(n14382), .Z(n11645) );
  COND11X1 U9012 ( .A(n15072), .B(n14389), .C(n14390), .D(n14877), .Z(n11646)
         );
  COND1XL U9013 ( .A(n14386), .B(n14385), .C(n15145), .Z(n11647) );
  CND4X1 U9014 ( .A(n14391), .B(n11645), .C(n11646), .D(n11647), .Z(n8729) );
  COND1XL U9015 ( .A(poly0_shifted[207]), .B(n18206), .C(n18163), .Z(n11648)
         );
  CND2X1 U9016 ( .A(n18119), .B(Poly0[207]), .Z(n11649) );
  COND1XL U9017 ( .A(n18119), .B(n11648), .C(n11649), .Z(n9370) );
  COND1XL U9018 ( .A(poly0_shifted[210]), .B(n18210), .C(n18172), .Z(n11650)
         );
  CND2X1 U9019 ( .A(n18119), .B(Poly0[210]), .Z(n11651) );
  COND1XL U9020 ( .A(n18119), .B(n11650), .C(n11651), .Z(n9367) );
  COND1XL U9021 ( .A(poly0_shifted[217]), .B(n18249), .C(n18196), .Z(n11652)
         );
  CND2X1 U9022 ( .A(n18119), .B(Poly0[217]), .Z(n11653) );
  COND1XL U9023 ( .A(n18119), .B(n11652), .C(n11653), .Z(n9360) );
  CMXI2X1 U9024 ( .A0(n14355), .A1(Poly8[90]), .S(Poly8[75]), .Z(n11654) );
  CND2X1 U9025 ( .A(n17156), .B(n11654), .Z(n11655) );
  CMXI2X1 U9026 ( .A0(n18249), .A1(Poly8[89]), .S(n17750), .Z(n11656) );
  CND2X1 U9027 ( .A(n11655), .B(n11656), .Z(n11312) );
  CANR2XL U9028 ( .A(n17652), .B(Poly12[124]), .C(poly12_shifted[124]), .D(
        n18017), .Z(n11657) );
  COND1XL U9029 ( .A(n17652), .B(n11978), .C(n11657), .Z(n10408) );
  CND2X1 U9030 ( .A(poly5_shifted[85]), .B(n17755), .Z(n11658) );
  CMXI2X1 U9031 ( .A0(Poly5[85]), .A1(n18241), .S(n17045), .Z(n11659) );
  CND2X1 U9032 ( .A(n11658), .B(n11659), .Z(n11441) );
  COND1XL U9033 ( .A(poly9_shifted[44]), .B(n13028), .C(n18153), .Z(n11660) );
  CND2X1 U9034 ( .A(n13351), .B(poly9_shifted[55]), .Z(n11661) );
  COND1XL U9035 ( .A(n13351), .B(n11660), .C(n11661), .Z(n11261) );
  COND1XL U9036 ( .A(poly0_shifted[212]), .B(n18082), .C(n18200), .Z(n11662)
         );
  CND2X1 U9037 ( .A(n18119), .B(Poly0[212]), .Z(n11663) );
  COND1XL U9038 ( .A(n18119), .B(n11662), .C(n11663), .Z(n9365) );
  COND1XL U9039 ( .A(poly0_shifted[197]), .B(n11988), .C(n18134), .Z(n11664)
         );
  CND2X1 U9040 ( .A(n18119), .B(poly0_shifted[215]), .Z(n11665) );
  COND1XL U9041 ( .A(n18119), .B(n11664), .C(n11665), .Z(n9380) );
  COND1XL U9042 ( .A(Poly10[40]), .B(Poly10[2]), .C(n18017), .Z(n11666) );
  CMXI2X1 U9043 ( .A0(n18160), .A1(Poly10[14]), .S(n17962), .Z(n11667) );
  COND4CX1 U9044 ( .A(Poly10[2]), .B(Poly10[40]), .C(n11666), .D(n11667), .Z(
        n11089) );
  CND2X1 U9045 ( .A(n12211), .B(poly2_shifted[23]), .Z(n11668) );
  COND4CX1 U9046 ( .A(n16753), .B(n16605), .C(n12211), .D(n11668), .Z(n8999)
         );
  COND1XL U9047 ( .A(n13522), .B(poly2_shifted[17]), .C(n18193), .Z(n11669) );
  CND2X1 U9048 ( .A(n12211), .B(poly2_shifted[29]), .Z(n11670) );
  COND1XL U9049 ( .A(n12211), .B(n11669), .C(n11670), .Z(n8993) );
  COND1XL U9050 ( .A(poly11_shifted[24]), .B(n13994), .C(n18091), .Z(n11671)
         );
  CND2X1 U9051 ( .A(n12185), .B(Poly11[24]), .Z(n11672) );
  COND1XL U9052 ( .A(n12185), .B(n11671), .C(n11672), .Z(n11165) );
  COND1XL U9053 ( .A(poly8_shifted[58]), .B(n18095), .C(n18094), .Z(n11673) );
  CND2X1 U9054 ( .A(n12287), .B(poly8_shifted[72]), .Z(n11674) );
  COND1XL U9055 ( .A(n12287), .B(n11673), .C(n11674), .Z(n11343) );
  CENX1 U9056 ( .A(dataselector[23]), .B(n17830), .Z(n11675) );
  CIVX1 U9057 ( .A(n17831), .Z(n11676) );
  CANR2X1 U9058 ( .A(n17832), .B(n18105), .C(dataselector[30]), .D(n11676), 
        .Z(n11677) );
  COND1XL U9059 ( .A(n17959), .B(n11675), .C(n11677), .Z(n8765) );
  COND1XL U9060 ( .A(poly3_shifted[22]), .B(n14487), .C(n18088), .Z(n11678) );
  CND2X1 U9061 ( .A(n15737), .B(poly3_shifted[36]), .Z(n11679) );
  COND1XL U9062 ( .A(n15737), .B(n11678), .C(n11679), .Z(n8918) );
  CND2X1 U9063 ( .A(poly5_shifted[77]), .B(n17238), .Z(n11680) );
  CMXI2X1 U9064 ( .A0(Poly5[77]), .A1(n18219), .S(n17045), .Z(n11681) );
  CND2X1 U9065 ( .A(n11680), .B(n11681), .Z(n11449) );
  CMXI2X1 U9066 ( .A0(n18099), .A1(poly10_shifted[39]), .S(n17962), .Z(n11682)
         );
  COND1XL U9067 ( .A(n15951), .B(Poly10[15]), .C(n17466), .Z(n11683) );
  COND4CX1 U9068 ( .A(Poly10[15]), .B(n15951), .C(n11683), .D(n11682), .Z(
        n11076) );
  CIVX1 U9069 ( .A(n13251), .Z(n11684) );
  CENX1 U9070 ( .A(Poly3[79]), .B(Poly3[46]), .Z(n11685) );
  CANR1XL U9071 ( .A(n14516), .B(n11685), .C(n12007), .Z(n11686) );
  COND11X1 U9072 ( .A(n18208), .B(Poly3[46]), .C(n12614), .D(n11686), .Z(
        n11687) );
  CMXI2X1 U9073 ( .A0(poly3_shifted[74]), .A1(n11687), .S(n12616), .Z(n11688)
         );
  COND11X1 U9074 ( .A(Poly3[79]), .B(n12615), .C(n11684), .D(n11688), .Z(n8880) );
  CENX1 U9075 ( .A(Poly12[118]), .B(Poly12[59]), .Z(n11689) );
  CANR1XL U9076 ( .A(n17994), .B(n11689), .C(n16381), .Z(n11690) );
  CIVX1 U9077 ( .A(n11689), .Z(n11691) );
  CANR2X1 U9078 ( .A(n12161), .B(poly12_shifted[91]), .C(n11691), .D(n17995), 
        .Z(n11692) );
  COND1XL U9079 ( .A(n12161), .B(n11690), .C(n11692), .Z(n10457) );
  COND1XL U9080 ( .A(n18116), .B(poly0_shifted[70]), .C(n18117), .Z(n11693) );
  CND2X1 U9081 ( .A(n12291), .B(poly0_shifted[88]), .Z(n11694) );
  COND1XL U9082 ( .A(n12291), .B(n11693), .C(n11694), .Z(n9507) );
  CEOX1 U9083 ( .A(Poly15[14]), .B(Poly15[47]), .Z(n11695) );
  CMX2GX1 U9084 ( .GN(n18228), .A0(n18040), .A1(n13940), .S(n11695), .Z(n11696) );
  CND2X1 U9085 ( .A(n18044), .B(Poly15[29]), .Z(n11697) );
  COND1XL U9086 ( .A(n11696), .B(n18044), .C(n11697), .Z(n9608) );
  CND2X1 U9087 ( .A(poly5_shifted[65]), .B(n17398), .Z(n11698) );
  CMXI2X1 U9088 ( .A0(poly5_shifted[79]), .A1(n14716), .S(n17045), .Z(n11699)
         );
  CND2X1 U9089 ( .A(n11698), .B(n11699), .Z(n11461) );
  CND2X1 U9090 ( .A(poly5_shifted[46]), .B(n17063), .Z(n11700) );
  CMXI2X1 U9091 ( .A0(poly5_shifted[60]), .A1(n18160), .S(n12942), .Z(n11701)
         );
  CND2X1 U9092 ( .A(n11700), .B(n11701), .Z(n11480) );
  CANR2X1 U9093 ( .A(n12175), .B(Poly8[9]), .C(Poly8[91]), .D(n16947), .Z(
        n11702) );
  COND1XL U9094 ( .A(n12175), .B(n12002), .C(n11702), .Z(n11392) );
  COND1XL U9095 ( .A(Poly14[290]), .B(Poly14[198]), .C(n17655), .Z(n11703) );
  CMXI2X1 U9096 ( .A0(n18034), .A1(Poly14[214]), .S(n12202), .Z(n11704) );
  COND4CX1 U9097 ( .A(Poly14[198]), .B(Poly14[290]), .C(n11703), .D(n11704), 
        .Z(n10191) );
  CND2X1 U9098 ( .A(n15050), .B(n15051), .Z(n11705) );
  CANR1XL U9099 ( .A(n15053), .B(n15054), .C(n12055), .Z(n11706) );
  CNR2X1 U9100 ( .A(n11705), .B(n11706), .Z(n15055) );
  COND1XL U9101 ( .A(n15168), .B(n14908), .C(n15153), .Z(n11707) );
  CND2IX1 U9102 ( .B(n14645), .A(n11707), .Z(n14921) );
  CAN4X1 U9103 ( .A(n12472), .B(n14909), .C(n15024), .D(n15270), .Z(n12046) );
  COND1XL U9104 ( .A(n13958), .B(n14966), .C(n15251), .Z(n11708) );
  COND11X1 U9105 ( .A(n14696), .B(n14697), .C(n11708), .D(n12216), .Z(n14700)
         );
  CNR2IX1 U9106 ( .B(n17136), .A(Poly11[78]), .Z(n14300) );
  CND2IX1 U9107 ( .B(n17628), .A(n16326), .Z(n15246) );
  CNR2IX1 U9108 ( .B(n18017), .A(Poly1[339]), .Z(n13362) );
  CNR2IXL U9109 ( .B(n18017), .A(Poly5[113]), .Z(n17940) );
  CND3XL U9110 ( .A(n17280), .B(Poly15[28]), .C(n16742), .Z(n13057) );
  CND2IX1 U9111 ( .B(Poly2[63]), .A(n17620), .Z(n12936) );
  CND2IX1 U9112 ( .B(Poly6[48]), .A(n17714), .Z(n13467) );
  COND1XL U9113 ( .A(Poly10[36]), .B(Poly10[41]), .C(n17714), .Z(n11709) );
  CANR1XL U9114 ( .A(Poly10[36]), .B(Poly10[41]), .C(n11709), .Z(n13572) );
  CNR2IX1 U9115 ( .B(n17714), .A(Poly12[120]), .Z(n14284) );
  CANR2X1 U9116 ( .A(n16877), .B(Poly7[25]), .C(n16839), .D(
        poly14_shifted[247]), .Z(n11710) );
  CANR2X1 U9117 ( .A(n16837), .B(poly14_shifted[68]), .C(poly13_shifted[457]), 
        .D(n12084), .Z(n11711) );
  CAN4X1 U9118 ( .A(n11710), .B(n11711), .C(n14527), .D(n14528), .Z(n14534) );
  CNR2X1 U9119 ( .A(n15318), .B(n15144), .Z(n11712) );
  CND3XL U9120 ( .A(n15142), .B(n15143), .C(n11712), .Z(n15146) );
  CIVX1 U9121 ( .A(n15247), .Z(n11713) );
  CND2X1 U9122 ( .A(n15248), .B(n17779), .Z(n11714) );
  CANR1XL U9123 ( .A(n15249), .B(n11713), .C(n11714), .Z(n15254) );
  CANR3X1 U9124 ( .A(n14889), .B(n12216), .C(n14885), .D(n14884), .Z(n11715)
         );
  CND3XL U9125 ( .A(n14898), .B(n14899), .C(n11715), .Z(n8719) );
  COND1XL U9126 ( .A(poly0_shifted[215]), .B(n11999), .C(n18203), .Z(n11716)
         );
  CND2X1 U9127 ( .A(n18119), .B(Poly0[215]), .Z(n11717) );
  COND1XL U9128 ( .A(n18119), .B(n11716), .C(n11717), .Z(n9362) );
  COND1XL U9129 ( .A(poly9_shifted[111]), .B(n18206), .C(n18163), .Z(n11718)
         );
  CND2X1 U9130 ( .A(n12262), .B(Poly9[111]), .Z(n11719) );
  COND1XL U9131 ( .A(n12262), .B(n11718), .C(n11719), .Z(n11194) );
  COND1XL U9132 ( .A(poly0_shifted[203]), .B(n16381), .C(n18150), .Z(n11720)
         );
  CND2X1 U9133 ( .A(n18119), .B(Poly0[203]), .Z(n11721) );
  COND1XL U9134 ( .A(n18119), .B(n11720), .C(n11721), .Z(n9374) );
  CND2X1 U9135 ( .A(Poly6[14]), .B(n13498), .Z(n11722) );
  COND3X1 U9136 ( .A(Poly6[14]), .B(n13408), .C(n11722), .D(n17721), .Z(n11723) );
  CMX2X1 U9137 ( .A0(n11723), .A1(Poly6[24]), .S(n13840), .Z(n9669) );
  COND1XL U9138 ( .A(poly0_shifted[211]), .B(n18176), .C(n18175), .Z(n11724)
         );
  CND2X1 U9139 ( .A(n18119), .B(Poly0[211]), .Z(n11725) );
  COND1XL U9140 ( .A(n18119), .B(n11724), .C(n11725), .Z(n9366) );
  COND1XL U9141 ( .A(poly4_shifted[21]), .B(n18241), .C(n18085), .Z(n11726) );
  CND2X1 U9142 ( .A(n18230), .B(Poly4[21]), .Z(n11727) );
  COND1XL U9143 ( .A(n18230), .B(n11726), .C(n11727), .Z(n8835) );
  CND2X1 U9144 ( .A(Poly8[90]), .B(n17063), .Z(n11728) );
  CND2X1 U9145 ( .A(n12175), .B(Poly8[8]), .Z(n11729) );
  COND3X1 U9146 ( .A(n12175), .B(n17163), .C(n11729), .D(n11728), .Z(n11393)
         );
  COND1XL U9147 ( .A(poly4_shifted[25]), .B(n18249), .C(n18196), .Z(n11730) );
  CND2X1 U9148 ( .A(n18230), .B(Poly4[25]), .Z(n11731) );
  COND1XL U9149 ( .A(n18230), .B(n11730), .C(n11731), .Z(n8831) );
  CND2X1 U9150 ( .A(n17312), .B(n17313), .Z(n11732) );
  COND3X1 U9151 ( .A(n17311), .B(n17310), .C(n17309), .D(n11983), .Z(n11733)
         );
  CMXI2X1 U9152 ( .A0(Poly2[37]), .A1(n11733), .S(n12021), .Z(n11734) );
  CND2X1 U9153 ( .A(n11732), .B(n11734), .Z(n8973) );
  CND2X1 U9154 ( .A(poly5_shifted[80]), .B(n17144), .Z(n11735) );
  CMXI2X1 U9155 ( .A0(Poly5[80]), .A1(n18167), .S(n17045), .Z(n11736) );
  CND2X1 U9156 ( .A(n11735), .B(n11736), .Z(n11446) );
  CANR2X1 U9157 ( .A(poly13_shifted[72]), .B(n17348), .C(n17969), .D(
        poly13_shifted[86]), .Z(n11737) );
  COND1XL U9158 ( .A(n17969), .B(n17163), .C(n11737), .Z(n10988) );
  COND1XL U9159 ( .A(poly8_shifted[39]), .B(n18138), .C(n18137), .Z(n11738) );
  CND2X1 U9160 ( .A(n12287), .B(poly8_shifted[53]), .Z(n11739) );
  COND1XL U9161 ( .A(n12287), .B(n11738), .C(n11739), .Z(n11362) );
  COND1XL U9162 ( .A(poly0_shifted[194]), .B(n12415), .C(n18126), .Z(n11740)
         );
  CND2X1 U9163 ( .A(n18119), .B(poly0_shifted[212]), .Z(n11741) );
  COND1XL U9164 ( .A(n18119), .B(n11740), .C(n11741), .Z(n9383) );
  COND1XL U9165 ( .A(poly8_shifted[44]), .B(n13028), .C(n18153), .Z(n11742) );
  CND2X1 U9166 ( .A(n12287), .B(poly8_shifted[58]), .Z(n11743) );
  COND1XL U9167 ( .A(n12287), .B(n11742), .C(n11743), .Z(n11357) );
  CND2X1 U9168 ( .A(n17962), .B(Poly10[2]), .Z(n11744) );
  COND4CX1 U9169 ( .A(n13756), .B(n16303), .C(n17962), .D(n11744), .Z(n11101)
         );
  CANR2X1 U9170 ( .A(n14448), .B(n13781), .C(dataselector[38]), .D(n16350), 
        .Z(n11745) );
  COND1XL U9171 ( .A(n14448), .B(n13780), .C(n17757), .Z(n11746) );
  CND2X1 U9172 ( .A(n11746), .B(n18252), .Z(n11747) );
  CND2X1 U9173 ( .A(n11745), .B(n11747), .Z(n8757) );
  CANR2X1 U9174 ( .A(n17314), .B(Poly0[162]), .C(poly0_shifted[162]), .D(
        n17215), .Z(n11748) );
  COND1XL U9175 ( .A(n17316), .B(n16303), .C(n11748), .Z(n9415) );
  CANR2X1 U9176 ( .A(n12170), .B(Poly7[55]), .C(poly7_shifted[55]), .D(n16326), 
        .Z(n11749) );
  COND1XL U9177 ( .A(n12170), .B(n12296), .C(n11749), .Z(n10049) );
  CANR2XL U9178 ( .A(n12161), .B(Poly12[92]), .C(poly12_shifted[92]), .D(
        n18017), .Z(n11750) );
  COND1XL U9179 ( .A(n12161), .B(n11978), .C(n11750), .Z(n10440) );
  CENX1 U9180 ( .A(Poly12[112]), .B(Poly12[23]), .Z(n11751) );
  CANR1XL U9181 ( .A(n17994), .B(n11751), .C(n18138), .Z(n11752) );
  CIVX1 U9182 ( .A(n11751), .Z(n11753) );
  CANR2X1 U9183 ( .A(n12598), .B(poly12_shifted[55]), .C(n11753), .D(n17995), 
        .Z(n11754) );
  COND1XL U9184 ( .A(n12598), .B(n11752), .C(n11754), .Z(n10493) );
  COND1XL U9185 ( .A(n18116), .B(Poly1[342]), .C(n18117), .Z(n11755) );
  CND2X1 U9186 ( .A(n18180), .B(poly1_shifted[17]), .Z(n11756) );
  COND1XL U9187 ( .A(n18180), .B(n11755), .C(n11756), .Z(n9351) );
  COND1XL U9188 ( .A(poly1_shifted[30]), .B(n18105), .C(n18104), .Z(n11757) );
  CND2X1 U9189 ( .A(n18180), .B(Poly1[30]), .Z(n11758) );
  COND1XL U9190 ( .A(n18180), .B(n11757), .C(n11758), .Z(n9327) );
  COND1XL U9191 ( .A(poly1_shifted[24]), .B(n13994), .C(n18091), .Z(n11759) );
  CND2X1 U9192 ( .A(n18180), .B(Poly1[24]), .Z(n11760) );
  COND1XL U9193 ( .A(n18180), .B(n11759), .C(n11760), .Z(n9333) );
  COND1XL U9194 ( .A(poly1_shifted[26]), .B(n18095), .C(n18094), .Z(n11761) );
  CND2X1 U9195 ( .A(n18180), .B(Poly1[26]), .Z(n11762) );
  COND1XL U9196 ( .A(n18180), .B(n11761), .C(n11762), .Z(n9331) );
  COND1XL U9197 ( .A(poly1_shifted[27]), .B(n18099), .C(n18098), .Z(n11763) );
  CND2X1 U9198 ( .A(n18180), .B(Poly1[27]), .Z(n11764) );
  COND1XL U9199 ( .A(n18180), .B(n11763), .C(n11764), .Z(n9330) );
  COND1XL U9200 ( .A(poly1_shifted[22]), .B(n14487), .C(n18088), .Z(n11765) );
  CND2X1 U9201 ( .A(n18180), .B(Poly1[22]), .Z(n11766) );
  COND1XL U9202 ( .A(n18180), .B(n11765), .C(n11766), .Z(n9335) );
  CND2XL U9203 ( .A(poly5_shifted[81]), .B(n18017), .Z(n11767) );
  CMXI2X1 U9204 ( .A0(Poly5[81]), .A1(n13522), .S(n17045), .Z(n11768) );
  CND2X1 U9205 ( .A(n11767), .B(n11768), .Z(n11445) );
  CENX1 U9206 ( .A(dataselector[10]), .B(n17828), .Z(n11769) );
  CIVX1 U9207 ( .A(n17831), .Z(n11770) );
  CANR2X1 U9208 ( .A(n17832), .B(n14297), .C(dataselector[17]), .D(n11770), 
        .Z(n11771) );
  COND1XL U9209 ( .A(n17829), .B(n11769), .C(n11771), .Z(n8778) );
  CND2X1 U9210 ( .A(Poly5[115]), .B(n17288), .Z(n11772) );
  CMXI2X1 U9211 ( .A0(Poly5[4]), .A1(n12004), .S(n17016), .Z(n11773) );
  CND2X1 U9212 ( .A(n11772), .B(n11773), .Z(n11522) );
  CANR2XL U9213 ( .A(n12299), .B(poly1_shifted[58]), .C(poly1_shifted[47]), 
        .D(n18017), .Z(n11774) );
  COND1XL U9214 ( .A(n12299), .B(n17196), .C(n11774), .Z(n9310) );
  CANR2X1 U9215 ( .A(n13040), .B(poly7_shifted[339]), .C(poly7_shifted[327]), 
        .D(n17206), .Z(n11775) );
  COND1XL U9216 ( .A(n13040), .B(n17718), .C(n11775), .Z(n9777) );
  COAN1X1 U9217 ( .A(Poly5[90]), .B(n13417), .C(n17163), .Z(n11776) );
  CND3XL U9218 ( .A(Poly5[90]), .B(n16326), .C(n12627), .Z(n11777) );
  CND2X1 U9219 ( .A(n12016), .B(poly5_shifted[118]), .Z(n11778) );
  COND3X1 U9220 ( .A(n13904), .B(n11776), .C(n11777), .D(n11778), .Z(n11422)
         );
  CND2X1 U9221 ( .A(poly5_shifted[48]), .B(n16479), .Z(n11779) );
  CMXI2X1 U9222 ( .A0(poly5_shifted[62]), .A1(n18167), .S(n12942), .Z(n11780)
         );
  CND2X1 U9223 ( .A(n11779), .B(n11780), .Z(n11478) );
  CND2X1 U9224 ( .A(poly5_shifted[69]), .B(n17538), .Z(n11781) );
  CMXI2X1 U9225 ( .A0(poly5_shifted[83]), .A1(n11990), .S(n17045), .Z(n11782)
         );
  CND2X1 U9226 ( .A(n11781), .B(n11782), .Z(n11457) );
  COND1XL U9227 ( .A(Poly14[297]), .B(Poly14[177]), .C(n17545), .Z(n11783) );
  CMXI2X1 U9228 ( .A0(n14361), .A1(Poly14[193]), .S(n12202), .Z(n11784) );
  COND4CX1 U9229 ( .A(Poly14[177]), .B(Poly14[297]), .C(n11783), .D(n11784), 
        .Z(n10212) );
  CANR2X1 U9230 ( .A(poly0_shifted[58]), .B(n17500), .C(n14159), .D(n18142), 
        .Z(n11785) );
  CENX1 U9231 ( .A(Poly0[22]), .B(Poly0[219]), .Z(n11786) );
  COND1XL U9232 ( .A(n17160), .B(n11786), .C(n11785), .Z(n9537) );
  CMXI2X1 U9233 ( .A0(n12199), .A1(Poly12[123]), .S(Poly12[93]), .Z(n11787) );
  CND2X1 U9234 ( .A(n17398), .B(n11787), .Z(n11788) );
  CMXI2X1 U9235 ( .A0(poly12_shifted[125]), .A1(n18219), .S(n18001), .Z(n11789) );
  CND2X1 U9236 ( .A(n11788), .B(n11789), .Z(n10423) );
  COND1XL U9237 ( .A(Poly7[234]), .B(Poly7[400]), .C(n17449), .Z(n11790) );
  CMXI2X1 U9238 ( .A0(n18034), .A1(poly7_shifted[258]), .S(n17574), .Z(n11791)
         );
  COND4CX1 U9239 ( .A(Poly7[400]), .B(Poly7[234]), .C(n11790), .D(n11791), .Z(
        n9858) );
  CMXI2X1 U9240 ( .A0(n13986), .A1(Poly13[527]), .S(Poly13[282]), .Z(n11792)
         );
  CND2X1 U9241 ( .A(n17642), .B(n11792), .Z(n11793) );
  CMXI2X1 U9242 ( .A0(n18142), .A1(poly13_shifted[310]), .S(n17615), .Z(n11794) );
  CND2X1 U9243 ( .A(n11793), .B(n11794), .Z(n10764) );
  CIVX1 U9244 ( .A(n17799), .Z(n11795) );
  CANR3X1 U9245 ( .A(datain[1]), .B(n11795), .C(n15159), .D(n14982), .Z(n14470) );
  CND2IX1 U9246 ( .B(Poly15[59]), .A(n17634), .Z(n16558) );
  CND2IX1 U9247 ( .B(n15153), .A(n17804), .Z(n15154) );
  CND4X1 U9248 ( .A(n14684), .B(n15260), .C(n12050), .D(n14558), .Z(n11796) );
  CND2X1 U9249 ( .A(n12216), .B(n11796), .Z(n12057) );
  CNR2IX1 U9250 ( .B(datain[4]), .A(n14967), .Z(n17768) );
  CND2IX1 U9251 ( .B(n14390), .A(n14912), .Z(n12460) );
  CEOX1 U9252 ( .A(Poly4[53]), .B(Poly4[57]), .Z(n13928) );
  CEOX1 U9253 ( .A(n17884), .B(scrambler[16]), .Z(n17854) );
  CND2IX1 U9254 ( .B(n14647), .A(n11969), .Z(n15093) );
  CND2IX1 U9255 ( .B(Poly6[53]), .A(n17705), .Z(n13452) );
  CANR2X1 U9256 ( .A(entrophy[6]), .B(n11974), .C(entrophy[12]), .D(n13945), 
        .Z(n11797) );
  CANR11X1 U9257 ( .A(n11797), .B(n13946), .C(n14965), .D(n15170), .Z(n11798)
         );
  CNR2X1 U9258 ( .A(n13954), .B(n15236), .Z(n11799) );
  CNR2X1 U9259 ( .A(n11798), .B(n11799), .Z(n13976) );
  CND2IX1 U9260 ( .B(Poly0[9]), .A(n12765), .Z(n12676) );
  CNR2IX1 U9261 ( .B(n18017), .A(Poly6[51]), .Z(n14005) );
  CNR2IX1 U9262 ( .B(n17705), .A(Poly6[47]), .Z(n13861) );
  CNR2IX1 U9263 ( .B(n17705), .A(Poly12[118]), .Z(n14107) );
  CNR2IX1 U9264 ( .B(n17238), .A(Poly12[113]), .Z(n14292) );
  CND2IX1 U9265 ( .B(n15145), .A(n12561), .Z(n12562) );
  CIVX1 U9266 ( .A(n15286), .Z(n11800) );
  CND4X1 U9267 ( .A(n15287), .B(n17765), .C(n15344), .D(n11800), .Z(n15289) );
  COND1XL U9268 ( .A(poly0_shifted[204]), .B(n13028), .C(n18153), .Z(n11801)
         );
  CND2X1 U9269 ( .A(n18119), .B(Poly0[204]), .Z(n11802) );
  COND1XL U9270 ( .A(n18119), .B(n11801), .C(n11802), .Z(n9373) );
  COND1XL U9271 ( .A(poly0_shifted[202]), .B(n12013), .C(n18147), .Z(n11803)
         );
  CND2X1 U9272 ( .A(n18119), .B(Poly0[202]), .Z(n11804) );
  COND1XL U9273 ( .A(n18119), .B(n11803), .C(n11804), .Z(n9375) );
  CENX1 U9274 ( .A(Poly11[57]), .B(Poly11[78]), .Z(n11805) );
  CMXI2X1 U9275 ( .A0(n18142), .A1(Poly11[72]), .S(n15843), .Z(n11806) );
  COND1XL U9276 ( .A(n17495), .B(n11805), .C(n11806), .Z(n11117) );
  COND1XL U9277 ( .A(poly0_shifted[199]), .B(n18138), .C(n18137), .Z(n11807)
         );
  CND2X1 U9278 ( .A(n18119), .B(poly0_shifted[217]), .Z(n11808) );
  COND1XL U9279 ( .A(n18119), .B(n11807), .C(n11808), .Z(n9378) );
  COND1XL U9280 ( .A(Poly12[116]), .B(n13602), .C(n17449), .Z(n11809) );
  CMXI2X1 U9281 ( .A0(n16381), .A1(poly12_shifted[59]), .S(n12598), .Z(n11810)
         );
  COND4CX1 U9282 ( .A(n13602), .B(Poly12[116]), .C(n11809), .D(n11810), .Z(
        n10489) );
  CND2X1 U9283 ( .A(n16960), .B(n16961), .Z(n11811) );
  CND2X1 U9284 ( .A(Poly6[18]), .B(n16956), .Z(n11812) );
  CND2X1 U9285 ( .A(n11812), .B(n16958), .Z(n11813) );
  COND3X1 U9286 ( .A(n11812), .B(n16959), .C(n11813), .D(n11978), .Z(n11814)
         );
  CMXI2X1 U9287 ( .A0(Poly6[28]), .A1(n11814), .S(n16962), .Z(n11815) );
  CND2X1 U9288 ( .A(n11811), .B(n11815), .Z(n9665) );
  COND1XL U9289 ( .A(poly12_shifted[16]), .B(n18167), .C(n18166), .Z(n11816)
         );
  CND2X1 U9290 ( .A(n12997), .B(Poly12[16]), .Z(n11817) );
  COND1XL U9291 ( .A(n12997), .B(n11816), .C(n11817), .Z(n10516) );
  CANR2X1 U9292 ( .A(n18198), .B(poly1_shifted[311]), .C(poly1_shifted[300]), 
        .D(n16326), .Z(n11818) );
  COND1XL U9293 ( .A(n18198), .B(n17087), .C(n11818), .Z(n9057) );
  COND1XL U9294 ( .A(poly1_shifted[23]), .B(n11999), .C(n18203), .Z(n11819) );
  CND2X1 U9295 ( .A(n18180), .B(Poly1[23]), .Z(n11820) );
  COND1XL U9296 ( .A(n18180), .B(n11819), .C(n11820), .Z(n9334) );
  COND1XL U9297 ( .A(poly0_shifted[200]), .B(n18142), .C(n18141), .Z(n11821)
         );
  CND2X1 U9298 ( .A(n18119), .B(poly0_shifted[218]), .Z(n11822) );
  COND1XL U9299 ( .A(n18119), .B(n11821), .C(n11822), .Z(n9377) );
  COND1XL U9300 ( .A(n13522), .B(poly9_shifted[49]), .C(n18193), .Z(n11823) );
  CND2X1 U9301 ( .A(n13351), .B(poly9_shifted[60]), .Z(n11824) );
  COND1XL U9302 ( .A(n13351), .B(n11823), .C(n11824), .Z(n11256) );
  CND2X1 U9303 ( .A(poly5_shifted[68]), .B(n17238), .Z(n11825) );
  CMXI2X1 U9304 ( .A0(poly5_shifted[82]), .A1(n12004), .S(n17045), .Z(n11826)
         );
  CND2X1 U9305 ( .A(n11825), .B(n11826), .Z(n11458) );
  CND2X1 U9306 ( .A(poly5_shifted[20]), .B(n17238), .Z(n11827) );
  CMXI2X1 U9307 ( .A0(poly5_shifted[34]), .A1(n18082), .S(n17016), .Z(n11828)
         );
  CND2X1 U9308 ( .A(n11827), .B(n11828), .Z(n11506) );
  COND1XL U9309 ( .A(poly9_shifted[89]), .B(n18249), .C(n18196), .Z(n11829) );
  CND2X1 U9310 ( .A(n17955), .B(Poly9[89]), .Z(n11830) );
  COND1XL U9311 ( .A(n17955), .B(n11829), .C(n11830), .Z(n11216) );
  CND3XL U9312 ( .A(Poly5[77]), .B(n17136), .C(n12627), .Z(n11831) );
  COND1XL U9313 ( .A(n13417), .B(Poly5[77]), .C(n17741), .Z(n11832) );
  CMXI2X1 U9314 ( .A0(n11832), .A1(Poly5[91]), .S(n17942), .Z(n11833) );
  CND2X1 U9315 ( .A(n11831), .B(n11833), .Z(n11435) );
  CENX1 U9316 ( .A(n15981), .B(dataselector[42]), .Z(n11834) );
  CIVX1 U9317 ( .A(n18252), .Z(n11835) );
  CANR2X1 U9318 ( .A(n17705), .B(n11834), .C(dataselector[49]), .D(n11835), 
        .Z(n11836) );
  COND1XL U9319 ( .A(n16139), .B(n17076), .C(n11836), .Z(n8746) );
  CND2X1 U9320 ( .A(poly5_shifted[79]), .B(n17705), .Z(n11837) );
  CMXI2X1 U9321 ( .A0(Poly5[79]), .A1(n18206), .S(n17045), .Z(n11838) );
  CND2X1 U9322 ( .A(n11837), .B(n11838), .Z(n11447) );
  CMXI2X1 U9323 ( .A0(n12013), .A1(Poly10[10]), .S(n17962), .Z(n11839) );
  CND2IX1 U9324 ( .B(n13572), .A(n11839), .Z(n11093) );
  CMXI2X1 U9325 ( .A0(n14355), .A1(Poly8[90]), .S(n13871), .Z(n11840) );
  CND2X1 U9326 ( .A(n17523), .B(n11840), .Z(n11841) );
  CMXI2X1 U9327 ( .A0(n18249), .A1(poly8_shifted[39]), .S(n12175), .Z(n11842)
         );
  CND2X1 U9328 ( .A(n11841), .B(n11842), .Z(n11376) );
  COND1XL U9329 ( .A(Poly15[57]), .B(Poly15[31]), .C(n16488), .Z(n11843) );
  CMXI2X1 U9330 ( .A0(n18160), .A1(Poly15[46]), .S(n17376), .Z(n11844) );
  COND4CX1 U9331 ( .A(Poly15[31]), .B(Poly15[57]), .C(n11843), .D(n11844), .Z(
        n9591) );
  CND2X1 U9332 ( .A(n12185), .B(poly11_shifted[23]), .Z(n11845) );
  COND3X1 U9333 ( .A(n12185), .B(n17163), .C(n11845), .D(n14190), .Z(n11181)
         );
  CNR2IX1 U9334 ( .B(Poly9[113]), .A(n15648), .Z(n11846) );
  CANR1XL U9335 ( .A(n17731), .B(poly9_shifted[19]), .C(n11846), .Z(n11847) );
  COND1XL U9336 ( .A(n17163), .B(n17731), .C(n11847), .Z(n11297) );
  CEOX1 U9337 ( .A(Poly2[28]), .B(Poly2[68]), .Z(n11848) );
  CENX1 U9338 ( .A(Poly2[64]), .B(n11848), .Z(n11849) );
  CNR2X1 U9339 ( .A(n17826), .B(n11849), .Z(n11850) );
  CANR1XL U9340 ( .A(n17306), .B(Poly2[40]), .C(n11850), .Z(n11851) );
  COND1XL U9341 ( .A(n17163), .B(n17306), .C(n11851), .Z(n8970) );
  COND1XL U9342 ( .A(n18116), .B(poly0_shifted[198]), .C(n18117), .Z(n11852)
         );
  CND2X1 U9343 ( .A(n18119), .B(poly0_shifted[216]), .Z(n11853) );
  COND1XL U9344 ( .A(n18119), .B(n11852), .C(n11853), .Z(n9379) );
  COND1XL U9345 ( .A(poly3_shifted[36]), .B(n12004), .C(n18131), .Z(n11854) );
  CND2X1 U9346 ( .A(n17262), .B(Poly3[36]), .Z(n11855) );
  COND1XL U9347 ( .A(n17262), .B(n11854), .C(n11855), .Z(n8904) );
  COND1XL U9348 ( .A(poly1_shifted[160]), .B(n12010), .C(n18185), .Z(n11856)
         );
  CND2X1 U9349 ( .A(n12210), .B(Poly1[160]), .Z(n11857) );
  COND1XL U9350 ( .A(n12210), .B(n11856), .C(n11857), .Z(n9197) );
  COND1XL U9351 ( .A(poly1_shifted[28]), .B(n12007), .C(n18224), .Z(n11858) );
  CND2X1 U9352 ( .A(n18180), .B(Poly1[28]), .Z(n11859) );
  COND1XL U9353 ( .A(n18180), .B(n11858), .C(n11859), .Z(n9329) );
  COND1XL U9354 ( .A(poly1_shifted[29]), .B(n18228), .C(n18227), .Z(n11860) );
  CND2X1 U9355 ( .A(n18180), .B(Poly1[29]), .Z(n11861) );
  COND1XL U9356 ( .A(n18180), .B(n11860), .C(n11861), .Z(n9328) );
  COND1XL U9357 ( .A(poly1_shifted[21]), .B(n18241), .C(n18085), .Z(n11862) );
  CND2X1 U9358 ( .A(n18180), .B(Poly1[21]), .Z(n11863) );
  COND1XL U9359 ( .A(n18180), .B(n11862), .C(n11863), .Z(n9336) );
  CEOX1 U9360 ( .A(Poly15[47]), .B(n13419), .Z(n11864) );
  CMX2GX1 U9361 ( .GN(n18105), .A0(n14323), .A1(n13420), .S(n11864), .Z(n11865) );
  CND2X1 U9362 ( .A(n18044), .B(Poly15[30]), .Z(n11866) );
  COND1XL U9363 ( .A(n11865), .B(n18044), .C(n11866), .Z(n9607) );
  COND1XL U9364 ( .A(poly7_shifted[58]), .B(n18095), .C(n18094), .Z(n11867) );
  CND2X1 U9365 ( .A(n12170), .B(Poly7[58]), .Z(n11868) );
  COND1XL U9366 ( .A(n12170), .B(n11867), .C(n11868), .Z(n10046) );
  COND1XL U9367 ( .A(poly7_shifted[52]), .B(n18082), .C(n18200), .Z(n11869) );
  CND2X1 U9368 ( .A(n12170), .B(Poly7[52]), .Z(n11870) );
  COND1XL U9369 ( .A(n12170), .B(n11869), .C(n11870), .Z(n10052) );
  COND1XL U9370 ( .A(poly14_shifted[178]), .B(n18210), .C(n18172), .Z(n11871)
         );
  CND2X1 U9371 ( .A(n13129), .B(Poly14[178]), .Z(n11872) );
  COND1XL U9372 ( .A(n13129), .B(n11871), .C(n11872), .Z(n10227) );
  COND1XL U9373 ( .A(poly14_shifted[169]), .B(n18189), .C(n18188), .Z(n11873)
         );
  CND2X1 U9374 ( .A(n13129), .B(Poly14[169]), .Z(n11874) );
  COND1XL U9375 ( .A(n13129), .B(n11873), .C(n11874), .Z(n10236) );
  COND1XL U9376 ( .A(poly9_shifted[14]), .B(n18160), .C(n18159), .Z(n11875) );
  CND2X1 U9377 ( .A(n17731), .B(Poly9[14]), .Z(n11876) );
  COND1XL U9378 ( .A(n17731), .B(n11875), .C(n11876), .Z(n11291) );
  COND1XL U9379 ( .A(poly5_shifted[88]), .B(n13994), .C(n18091), .Z(n11877) );
  CND2X1 U9380 ( .A(n17942), .B(Poly5[88]), .Z(n11878) );
  COND1XL U9381 ( .A(n17942), .B(n11877), .C(n11878), .Z(n11438) );
  CND2X1 U9382 ( .A(poly5_shifted[87]), .B(n18234), .Z(n11879) );
  CMXI2X1 U9383 ( .A0(Poly5[87]), .A1(n11999), .S(n17045), .Z(n11880) );
  CND2X1 U9384 ( .A(n11879), .B(n11880), .Z(n11439) );
  CND2X1 U9385 ( .A(poly5_shifted[76]), .B(n17535), .Z(n11881) );
  CMXI2X1 U9386 ( .A0(Poly5[76]), .A1(n13028), .S(n17045), .Z(n11882) );
  CND2X1 U9387 ( .A(n11881), .B(n11882), .Z(n11450) );
  CND2X1 U9388 ( .A(poly5_shifted[83]), .B(n17285), .Z(n11883) );
  CMXI2X1 U9389 ( .A0(Poly5[83]), .A1(n18176), .S(n17045), .Z(n11884) );
  CND2X1 U9390 ( .A(n11883), .B(n11884), .Z(n11443) );
  CANR2X1 U9391 ( .A(n18191), .B(poly1_shifted[278]), .C(poly1_shifted[267]), 
        .D(n17288), .Z(n11885) );
  COND1XL U9392 ( .A(n18191), .B(n16605), .C(n11885), .Z(n9090) );
  CANR2X1 U9393 ( .A(n18198), .B(poly1_shifted[301]), .C(poly1_shifted[290]), 
        .D(n16326), .Z(n11886) );
  COND1XL U9394 ( .A(n18198), .B(n16775), .C(n11886), .Z(n9067) );
  CANR2X1 U9395 ( .A(n17217), .B(poly7_shifted[127]), .C(poly7_shifted[115]), 
        .D(n16326), .Z(n11887) );
  COND1XL U9396 ( .A(n17217), .B(n17658), .C(n11887), .Z(n9989) );
  CND2X1 U9397 ( .A(poly5_shifted[75]), .B(n18234), .Z(n11888) );
  CMXI2X1 U9398 ( .A0(poly5_shifted[89]), .A1(n16381), .S(n17045), .Z(n11889)
         );
  CND2X1 U9399 ( .A(n11888), .B(n11889), .Z(n11451) );
  CIVX1 U9400 ( .A(n16565), .Z(n11890) );
  CANR1XL U9401 ( .A(n11890), .B(poly15_shifted[58]), .C(n13056), .Z(n11891)
         );
  CND2X1 U9402 ( .A(n13057), .B(n11891), .Z(n9594) );
  CND2X1 U9403 ( .A(poly5_shifted[71]), .B(n17362), .Z(n11892) );
  CMXI2X1 U9404 ( .A0(poly5_shifted[85]), .A1(n18138), .S(n17045), .Z(n11893)
         );
  CND2X1 U9405 ( .A(n11892), .B(n11893), .Z(n11455) );
  CND2X1 U9406 ( .A(poly5_shifted[67]), .B(n17535), .Z(n11894) );
  CMXI2X1 U9407 ( .A0(poly5_shifted[81]), .A1(n18053), .S(n17045), .Z(n11895)
         );
  CND2X1 U9408 ( .A(n11894), .B(n11895), .Z(n11459) );
  CND2X1 U9409 ( .A(poly5_shifted[72]), .B(n16427), .Z(n11896) );
  CMXI2X1 U9410 ( .A0(poly5_shifted[86]), .A1(n18142), .S(n17045), .Z(n11897)
         );
  CND2X1 U9411 ( .A(n11896), .B(n11897), .Z(n11454) );
  CMX2GX1 U9412 ( .GN(n18167), .A0(n17368), .A1(n12936), .S(Poly2[36]), .Z(
        n11898) );
  CND2X1 U9413 ( .A(n17306), .B(Poly2[48]), .Z(n11899) );
  COND1XL U9414 ( .A(n11898), .B(n17306), .C(n11899), .Z(n8962) );
  COND1XL U9415 ( .A(poly14_shifted[171]), .B(n16381), .C(n18150), .Z(n11900)
         );
  CND2X1 U9416 ( .A(n13129), .B(Poly14[171]), .Z(n11901) );
  COND1XL U9417 ( .A(n13129), .B(n11900), .C(n11901), .Z(n10234) );
  COND1XL U9418 ( .A(poly13_shifted[165]), .B(n11984), .C(n18134), .Z(n11902)
         );
  CND2X1 U9419 ( .A(n13014), .B(Poly13[165]), .Z(n11903) );
  COND1XL U9420 ( .A(n13014), .B(n11902), .C(n11903), .Z(n10895) );
  CIVX1 U9421 ( .A(n17831), .Z(n11904) );
  CANR2X1 U9422 ( .A(n17832), .B(n18138), .C(dataselector[7]), .D(n11904), .Z(
        n11905) );
  CENX1 U9423 ( .A(n17820), .B(dataselector[0]), .Z(n11906) );
  COND1XL U9424 ( .A(n17829), .B(n11906), .C(n11905), .Z(n8788) );
  CANR2X1 U9425 ( .A(Poly0[8]), .B(n17503), .C(Poly0[210]), .D(n17401), .Z(
        n11907) );
  COND1XL U9426 ( .A(n17506), .B(n17163), .C(n11907), .Z(n9569) );
  CMXI2X1 U9427 ( .A0(n14364), .A1(Poly1[345]), .S(Poly1[62]), .Z(n11908) );
  CND2X1 U9428 ( .A(n17121), .B(n11908), .Z(n11909) );
  CMXI2X1 U9429 ( .A0(n18189), .A1(poly1_shifted[84]), .S(n12012), .Z(n11910)
         );
  CND2X1 U9430 ( .A(n11909), .B(n11910), .Z(n9284) );
  CMXI2X1 U9431 ( .A0(n14360), .A1(Poly13[520]), .S(Poly13[275]), .Z(n11911)
         );
  CND2X1 U9432 ( .A(n16985), .B(n11911), .Z(n11912) );
  CMXI2X1 U9433 ( .A0(n14361), .A1(poly13_shifted[303]), .S(n17615), .Z(n11913) );
  CND2X1 U9434 ( .A(n11912), .B(n11913), .Z(n10771) );
  CMXI2X1 U9435 ( .A0(n12784), .A1(Poly12[121]), .S(Poly12[91]), .Z(n11914) );
  CND2X1 U9436 ( .A(n16695), .B(n11914), .Z(n11915) );
  CMXI2X1 U9437 ( .A0(poly12_shifted[123]), .A1(n16381), .S(n18001), .Z(n11916) );
  CND2X1 U9438 ( .A(n11915), .B(n11916), .Z(n10425) );
  CMXI2X1 U9439 ( .A0(n13592), .A1(Poly1[344]), .S(Poly1[61]), .Z(n11917) );
  CND2X1 U9440 ( .A(n17375), .B(n11917), .Z(n11918) );
  CMXI2X1 U9441 ( .A0(n18142), .A1(poly1_shifted[83]), .S(n12012), .Z(n11919)
         );
  CND2X1 U9442 ( .A(n11918), .B(n11919), .Z(n9285) );
  CMXI2X1 U9443 ( .A0(n14356), .A1(Poly1[341]), .S(Poly1[58]), .Z(n11920) );
  CND2X1 U9444 ( .A(n17105), .B(n11920), .Z(n11921) );
  CMXI2X1 U9445 ( .A0(n11990), .A1(poly1_shifted[80]), .S(n12012), .Z(n11922)
         );
  CND2X1 U9446 ( .A(n11921), .B(n11922), .Z(n9288) );
  CMXI2X1 U9447 ( .A0(n12003), .A1(poly7_shifted[267]), .S(n17574), .Z(n11923)
         );
  COND1XL U9448 ( .A(Poly7[243]), .B(Poly7[409]), .C(n17348), .Z(n11924) );
  COND4CX1 U9449 ( .A(Poly7[409]), .B(Poly7[243]), .C(n11924), .D(n11923), .Z(
        n9849) );
  COND1XL U9450 ( .A(Poly14[287]), .B(Poly14[167]), .C(n17466), .Z(n11925) );
  CMXI2X1 U9451 ( .A0(n11999), .A1(poly14_shifted[199]), .S(n13129), .Z(n11926) );
  COND4CX1 U9452 ( .A(Poly14[167]), .B(Poly14[287]), .C(n11925), .D(n11926), 
        .Z(n10222) );
  COND1XL U9453 ( .A(Poly14[286]), .B(Poly14[166]), .C(n18047), .Z(n11927) );
  CMXI2X1 U9454 ( .A0(n18034), .A1(poly14_shifted[198]), .S(n13129), .Z(n11928) );
  COND4CX1 U9455 ( .A(Poly14[166]), .B(Poly14[286]), .C(n11927), .D(n11928), 
        .Z(n10223) );
  CMXI2X1 U9456 ( .A0(n14363), .A1(Poly13[521]), .S(Poly13[276]), .Z(n11929)
         );
  CND2X1 U9457 ( .A(n16307), .B(n11929), .Z(n11930) );
  CMXI2X1 U9458 ( .A0(n13428), .A1(poly13_shifted[304]), .S(n17615), .Z(n11931) );
  CND2X1 U9459 ( .A(n11930), .B(n11931), .Z(n10770) );
  CMXI2X1 U9460 ( .A0(n14362), .A1(Poly13[515]), .S(Poly13[388]), .Z(n11932)
         );
  CND2X1 U9461 ( .A(n17209), .B(n11932), .Z(n11933) );
  CMXI2X1 U9462 ( .A0(n18210), .A1(poly13_shifted[416]), .S(n17043), .Z(n11934) );
  CND2X1 U9463 ( .A(n11933), .B(n11934), .Z(n10658) );
  CENX1 U9464 ( .A(Poly13[168]), .B(Poly13[527]), .Z(n11935) );
  CMXI2X1 U9465 ( .A0(n14487), .A1(poly13_shifted[196]), .S(n13014), .Z(n11936) );
  COND1XL U9466 ( .A(n17160), .B(n11935), .C(n11936), .Z(n10878) );
  CMXI2X1 U9467 ( .A0(n13591), .A1(Poly5[114]), .S(Poly5[92]), .Z(n11937) );
  CND2X1 U9468 ( .A(n17174), .B(n11937), .Z(n11938) );
  CMXI2X1 U9469 ( .A0(n12013), .A1(poly5_shifted[120]), .S(n15403), .Z(n11939)
         );
  CND2X1 U9470 ( .A(n11938), .B(n11939), .Z(n11420) );
  CENX1 U9471 ( .A(Poly2[33]), .B(n17692), .Z(n11940) );
  CND2X1 U9472 ( .A(n13553), .B(n11940), .Z(n11941) );
  COND1XL U9473 ( .A(n16753), .B(n11940), .C(n12949), .Z(n11942) );
  CMXI2X1 U9474 ( .A0(n11942), .A1(poly2_shifted[57]), .S(n17306), .Z(n11943)
         );
  CND2X1 U9475 ( .A(n11941), .B(n11943), .Z(n8965) );
  CEOX1 U9476 ( .A(Poly7[399]), .B(Poly7[19]), .Z(n11944) );
  CANR2X1 U9477 ( .A(n18018), .B(poly7_shifted[43]), .C(n11944), .D(n18017), 
        .Z(n11945) );
  COND1XL U9478 ( .A(n18019), .B(n18183), .C(n11945), .Z(n10073) );
  CANR2X1 U9479 ( .A(n12287), .B(poly8_shifted[46]), .C(poly8_shifted[32]), 
        .D(n18017), .Z(n11946) );
  COND1XL U9480 ( .A(n12287), .B(n17751), .C(n11946), .Z(n11369) );
  CENX1 U9481 ( .A(Poly12[120]), .B(Poly12[60]), .Z(n11947) );
  CANR1XL U9482 ( .A(n17994), .B(n11947), .C(n13028), .Z(n11948) );
  CIVX1 U9483 ( .A(n11947), .Z(n11949) );
  CANR2X1 U9484 ( .A(n12161), .B(poly12_shifted[92]), .C(n11949), .D(n17995), 
        .Z(n11950) );
  COND1XL U9485 ( .A(n12161), .B(n11948), .C(n11950), .Z(n10456) );
  CANR4CX1 U9486 ( .A(n15330), .B(n11971), .C(entrophy[3]), .D(n14544), .Z(
        n11951) );
  COND1XL U9487 ( .A(n14563), .B(n14562), .C(n15220), .Z(n11952) );
  CND4X1 U9488 ( .A(n14564), .B(n14565), .C(n11951), .D(n11952), .Z(n8701) );
  CANR2X1 U9489 ( .A(n18028), .B(poly7_shifted[327]), .C(poly7_shifted[315]), 
        .D(n18017), .Z(n11953) );
  COND1XL U9490 ( .A(n18028), .B(n17741), .C(n11953), .Z(n9789) );
  CMXI2X1 U9491 ( .A0(n14354), .A1(Poly10[35]), .S(Poly10[14]), .Z(n11954) );
  CND2X1 U9492 ( .A(n16427), .B(n11954), .Z(n11955) );
  CMXI2X1 U9493 ( .A0(n18095), .A1(Poly10[26]), .S(n17962), .Z(n11956) );
  CND2X1 U9494 ( .A(n11955), .B(n11956), .Z(n11077) );
  CMXI2X1 U9495 ( .A0(n18095), .A1(Poly9[26]), .S(n17731), .Z(n11957) );
  COND1XL U9496 ( .A(Poly9[107]), .B(Poly9[15]), .C(n17504), .Z(n11958) );
  COND4CX1 U9497 ( .A(Poly9[15]), .B(Poly9[107]), .C(n11958), .D(n11957), .Z(
        n11279) );
  CMXI2X1 U9498 ( .A0(n16381), .A1(Poly11[75]), .S(n15843), .Z(n11959) );
  CENX1 U9499 ( .A(Poly11[60]), .B(Poly11[81]), .Z(n11960) );
  COND1XL U9500 ( .A(n15673), .B(n11960), .C(n11959), .Z(n11114) );
  CAN4X1 U9501 ( .A(n16720), .B(n16721), .C(n16722), .D(n16723), .Z(n11961) );
  CND4X1 U9502 ( .A(n16736), .B(n16737), .C(n16738), .D(n11961), .Z(n11962) );
  CAOR2X1 U9503 ( .A(polydata[2]), .B(n17744), .C(n16886), .D(n11962), .Z(
        n8686) );
  COND2X1 U9504 ( .A(n15361), .B(n17090), .C(n17495), .D(n15418), .Z(n11963)
         );
  CAOR1X1 U9505 ( .A(n15378), .B(poly5_shifted[59]), .C(n11963), .Z(n11481) );
  CMXI2X1 U9506 ( .A0(n18099), .A1(Poly4[59]), .S(n12153), .Z(n11964) );
  CEOX1 U9507 ( .A(n13858), .B(n13857), .Z(n11965) );
  COND1XL U9508 ( .A(Poly4[51]), .B(n11965), .C(n17178), .Z(n11966) );
  COND4CX1 U9509 ( .A(n11965), .B(Poly4[51]), .C(n11966), .D(n11964), .Z(n8797) );
  CND2X2 U9510 ( .A(n12068), .B(dataselector[57]), .Z(n16349) );
  CND2X2 U9511 ( .A(n12068), .B(dataselector[5]), .Z(n12385) );
  CAN2X1 U9512 ( .A(n12068), .B(n13479), .Z(n13781) );
  CANR4CX2 U9513 ( .A(n16740), .B(n16743), .C(n12005), .D(n17376), .Z(n16741)
         );
  CND3X1 U9514 ( .A(n12496), .B(n12495), .C(n12494), .Z(n8703) );
  CIVX2 U9515 ( .A(n12173), .Z(n11967) );
  CAOR1X1 U9516 ( .A(n15309), .B(n14078), .C(n14077), .Z(n11968) );
  CNR2X2 U9517 ( .A(n11968), .B(n14076), .Z(n14101) );
  CIVDX2 U9518 ( .A(n17785), .Z0(n15309) );
  COND4CXL U9519 ( .A(n17779), .B(n14075), .C(n12055), .D(n14074), .Z(n14076)
         );
  CANR2XL U9520 ( .A(n12067), .B(poly12_shifted[126]), .C(n16872), .D(
        poly9_shifted[80]), .Z(n12078) );
  CANR2XL U9521 ( .A(n16863), .B(poly5_shifted[76]), .C(n16872), .D(Poly6[33]), 
        .Z(n12429) );
  CNR2X2 U9522 ( .A(n14788), .B(n14387), .Z(n14864) );
  CANR3X2 U9523 ( .A(n15314), .B(n14939), .C(n14938), .D(n14937), .Z(n14940)
         );
  COR2X1 U9524 ( .A(n17799), .B(n17798), .Z(n17802) );
  CND4X1 U9525 ( .A(n14989), .B(n14988), .C(n14987), .D(n14986), .Z(n14990) );
  CANR2X1 U9526 ( .A(n15034), .B(n14951), .C(scrambler[2]), .D(n17959), .Z(
        n14086) );
  COND1X4 U9527 ( .A(n12356), .B(n12404), .C(n17829), .Z(n13120) );
  COR2X1 U9528 ( .A(addr[3]), .B(addr[2]), .Z(n12356) );
  CNIVX12 U9529 ( .A(n12165), .Z(n17829) );
  CAOR1X1 U9530 ( .A(datain[3]), .B(n17812), .C(n14959), .Z(n14975) );
  CND2X2 U9531 ( .A(n15256), .B(dataselector[14]), .Z(n15168) );
  CIVDX3 U9532 ( .A(n12028), .Z0(n12173), .Z1(n12124) );
  CANR1X2 U9533 ( .A(n15145), .B(n14703), .C(n14702), .Z(n14710) );
  CND2X2 U9534 ( .A(n12704), .B(n13120), .Z(n17942) );
  CND2X1 U9535 ( .A(n12396), .B(n13120), .Z(n17411) );
  COND4CXL U9536 ( .A(entrophy[5]), .B(n15354), .C(n15353), .D(n14875), .Z(
        n15355) );
  CNR2X2 U9537 ( .A(addr[9]), .B(addr[11]), .Z(n12150) );
  CNR2X4 U9538 ( .A(n11973), .B(n15110), .Z(n14797) );
  CAN2X2 U9539 ( .A(n11969), .B(n17805), .Z(n11973) );
  CNIVX4 U9540 ( .A(pushin), .Z(n12028) );
  CIVDX2 U9541 ( .A(n13958), .Z0(n14680), .Z1(n14472) );
  CND3X2 U9542 ( .A(n12150), .B(n12149), .C(write), .Z(n12158) );
  CNR2X2 U9543 ( .A(addr[10]), .B(addr[8]), .Z(n12149) );
  COND1X1 U9544 ( .A(n16565), .B(n16564), .C(n16563), .Z(n9595) );
  CANR1X1 U9545 ( .A(n16562), .B(n16561), .C(n16560), .Z(n16563) );
  COND1X1 U9546 ( .A(n16565), .B(n14321), .C(n13022), .Z(n9589) );
  CANR1X1 U9547 ( .A(n16562), .B(Poly15[33]), .C(n13021), .Z(n13022) );
  CND2X2 U9548 ( .A(n12017), .B(n15583), .Z(n17430) );
  CIVX8 U9549 ( .A(n14454), .Z(n15218) );
  CIVDX2 U9550 ( .A(n12072), .Z0(n12064), .Z1(n12266) );
  CANR4CX2 U9551 ( .A(n15311), .B(n15310), .C(n15309), .D(n15308), .Z(n15317)
         );
  COND1X4 U9552 ( .A(n12261), .B(n12260), .C(n17495), .Z(n13189) );
  CIVX2 U9553 ( .A(n12031), .Z(n12072) );
  CNIVX4 U9554 ( .A(n14454), .Z(n15319) );
  CANR1X2 U9555 ( .A(n11977), .B(n12242), .C(n12068), .Z(n11976) );
  CIVX20 U9556 ( .A(n11976), .Z(n13267) );
  CIVX20 U9557 ( .A(n12261), .Z(n11977) );
  CNIVX12 U9558 ( .A(n12173), .Z(n17495) );
  CIVX3 U9559 ( .A(n14958), .Z(n15330) );
  CND2X2 U9560 ( .A(n12031), .B(dataselector[8]), .Z(n16249) );
  CIVDX3 U9561 ( .A(n12027), .Z0(n15145), .Z1(n17763) );
  CND2X2 U9562 ( .A(n17829), .B(lfsrdin[28]), .Z(n11978) );
  CND2X1 U9563 ( .A(n17829), .B(lfsrdin[28]), .Z(n18039) );
  CANR2X1 U9564 ( .A(entrophy[10]), .B(n17787), .C(n15314), .D(n15313), .Z(
        n15315) );
  CIVX8 U9565 ( .A(n17778), .Z(n12216) );
  CMXI2XL U9566 ( .A0(n12007), .A1(poly14_shifted[236]), .S(n12202), .Z(n14741) );
  CMXI2XL U9567 ( .A0(n12007), .A1(poly7_shifted[264]), .S(n17574), .Z(n14344)
         );
  CMXI2XL U9568 ( .A0(n12007), .A1(poly14_shifted[204]), .S(n13129), .Z(n14304) );
  CMXI2XL U9569 ( .A0(n12007), .A1(poly7_shifted[72]), .S(n12170), .Z(n13917)
         );
  CMXI2XL U9570 ( .A0(n12007), .A1(poly8_shifted[42]), .S(n12175), .Z(n13868)
         );
  CMXI2XL U9571 ( .A0(n12007), .A1(Poly8[92]), .S(n17750), .Z(n13827) );
  CMXI2XL U9572 ( .A0(n12007), .A1(poly13_shifted[298]), .S(n17592), .Z(n13821) );
  CMXI2XL U9573 ( .A0(n12007), .A1(poly10_shifted[40]), .S(n17962), .Z(n13732)
         );
  CMXI2XL U9574 ( .A0(n12007), .A1(poly13_shifted[426]), .S(n17043), .Z(n13566) );
  CMXI2XL U9575 ( .A0(n12007), .A1(Poly11[60]), .S(n17683), .Z(n13508) );
  CANR2XL U9576 ( .A(n15880), .B(poly0_shifted[142]), .C(n12007), .D(n16274), 
        .Z(n13696) );
  CIVX2 U9577 ( .A(n17732), .Z(n11979) );
  CIVX2 U9578 ( .A(n17732), .Z(n11980) );
  CIVDX1 U9579 ( .A(n11979), .Z0(n11981), .Z1(n11982) );
  CIVDX1 U9580 ( .A(n11979), .Z0(n11983), .Z1(n11984) );
  CIVDX1 U9581 ( .A(n11979), .Z0(n11985), .Z1(n11986) );
  CIVDX1 U9582 ( .A(n11979), .Z0(n11987), .Z1(n11988) );
  CIVDX1 U9583 ( .A(n11980), .Z0(n11989), .Z1(n11990) );
  CIVDX1 U9584 ( .A(n11980), .Z0(n11991), .Z1(n11992) );
  CIVDX1 U9585 ( .A(n11980), .Z0(n11993), .Z1(n11994) );
  CIVDX1 U9586 ( .A(n11980), .Z0(n11995), .Z1(n11996) );
  CND2X1 U9587 ( .A(n17495), .B(lfsrdin[5]), .Z(n17732) );
  CNIVX3 U9588 ( .A(n12024), .Z(n17160) );
  CIVX2 U9589 ( .A(n15648), .Z(n17634) );
  CND2X4 U9590 ( .A(n13267), .B(n12395), .Z(n17306) );
  CIVDX1 U9591 ( .A(n17306), .Z0(n12021), .Z1(n12022) );
  CIVDX4 U9592 ( .A(n18046), .Z0(n17376), .Z1(n16565) );
  CIVDX1 U9593 ( .A(n13421), .Z0(n11998), .Z1(n17747) );
  CND2X2 U9594 ( .A(n12704), .B(n13266), .Z(n15378) );
  CIVX3 U9595 ( .A(n12024), .Z(n12068) );
  CND2X1 U9596 ( .A(n17959), .B(lfsrdin[1]), .Z(n17711) );
  CNIVX12 U9597 ( .A(n12024), .Z(n15648) );
  CND2X2 U9598 ( .A(n12572), .B(lfsrdin[6]), .Z(n17757) );
  CIVDX2 U9599 ( .A(n16391), .Z0(n18082), .Z1(n17707) );
  CIVX3 U9600 ( .A(n17163), .Z(n18142) );
  CND2X4 U9601 ( .A(n17826), .B(lfsrdin[8]), .Z(n17163) );
  CNIVX4 U9602 ( .A(n12165), .Z(n15673) );
  CIVDX1 U9603 ( .A(n13354), .Z0(n12001), .Z1(n12002) );
  CND2X1 U9604 ( .A(n17744), .B(lfsrdin[9]), .Z(n13354) );
  CND2X1 U9605 ( .A(n17959), .B(lfsrdin[31]), .Z(n12968) );
  CIVDX3 U9606 ( .A(n12764), .Z0(n18160), .Z1(n17699) );
  CND2X1 U9607 ( .A(n17804), .B(dataselector[14]), .Z(n14963) );
  CND2X4 U9608 ( .A(n12017), .B(n13118), .Z(n13014) );
  CND2X4 U9609 ( .A(n12017), .B(n12991), .Z(n17491) );
  CND2X1 U9610 ( .A(n17959), .B(lfsrdin[12]), .Z(n17218) );
  CIVDX2 U9611 ( .A(n17218), .Z0(n13028), .Z1(n17087) );
  CND2X4 U9612 ( .A(n12017), .B(n13266), .Z(n17974) );
  CND2X4 U9613 ( .A(n12017), .B(n13145), .Z(n17982) );
  CND2X4 U9614 ( .A(n12017), .B(n12988), .Z(n17987) );
  CND2X4 U9615 ( .A(n12017), .B(n13128), .Z(n17667) );
  CND2X2 U9616 ( .A(n17495), .B(n14944), .Z(n17831) );
  CIVDX3 U9617 ( .A(n17831), .Z0(n16410), .Z1(n15799) );
  CIVDX2 U9618 ( .A(n12148), .Z0(n12004), .Z1(n12005) );
  CND2XL U9619 ( .A(n17829), .B(lfsrdin[4]), .Z(n12148) );
  CNR2X4 U9620 ( .A(n12115), .B(n12101), .Z(n12084) );
  CIVDX4 U9621 ( .A(n15042), .Z0(n17804), .Z1(n15334) );
  CNR2X4 U9622 ( .A(n12115), .B(n12112), .Z(n12067) );
  CIVDX1 U9623 ( .A(n12273), .Z0(n18241), .Z1(n17036) );
  CNIVX2 U9624 ( .A(n12572), .Z(n17259) );
  CIVDX1 U9625 ( .A(n13367), .Z1(n17735) );
  CIVDX1 U9626 ( .A(n13367), .Z0(n18095), .Z1(n17305) );
  CND2X1 U9627 ( .A(n17959), .B(lfsrdin[26]), .Z(n13367) );
  CIVDX2 U9628 ( .A(n17718), .Z0(n18138), .Z1(n16939) );
  CND2X2 U9629 ( .A(n17744), .B(lfsrdin[7]), .Z(n17718) );
  CIVDX4 U9630 ( .A(n14132), .Z0(n14695), .Z1(n14226) );
  CND2X4 U9631 ( .A(n17744), .B(lfsrdin[3]), .Z(n13275) );
  CIVX4 U9632 ( .A(n13275), .Z(n18053) );
  CND2X1 U9633 ( .A(n17495), .B(lfsrdin[2]), .Z(n16387) );
  CND2X4 U9634 ( .A(n13267), .B(n13145), .Z(n17332) );
  CND2X4 U9635 ( .A(n13100), .B(n13266), .Z(n17471) );
  CND2X4 U9636 ( .A(n12250), .B(n13145), .Z(n12153) );
  CND2X4 U9637 ( .A(n13100), .B(n12610), .Z(n17273) );
  CND2X1 U9638 ( .A(n12068), .B(n18257), .Z(n14852) );
  CND2X2 U9639 ( .A(n17959), .B(lfsrdin[30]), .Z(n13418) );
  CND2X4 U9640 ( .A(n13189), .B(n13093), .Z(n12262) );
  CND2X2 U9641 ( .A(n17744), .B(lfsrdin[22]), .Z(n17753) );
  CND2X4 U9642 ( .A(n13100), .B(n13118), .Z(n13070) );
  CND2X4 U9643 ( .A(n13100), .B(n13227), .Z(n12625) );
  CND2X4 U9644 ( .A(n13100), .B(n13093), .Z(n12206) );
  CND2X4 U9645 ( .A(n13100), .B(n13128), .Z(n12977) );
  CND2X4 U9646 ( .A(n12250), .B(n13120), .Z(n15737) );
  CND2X4 U9647 ( .A(n13100), .B(n13145), .Z(n13040) );
  CND2X4 U9648 ( .A(n12396), .B(n13093), .Z(n12185) );
  CND2X4 U9649 ( .A(n13878), .B(n13266), .Z(n12958) );
  CND2X4 U9650 ( .A(n13267), .B(n12988), .Z(n12211) );
  CND2X4 U9651 ( .A(n13189), .B(n13877), .Z(n12287) );
  CND2X4 U9652 ( .A(n13123), .B(n12994), .Z(n12900) );
  CND2X4 U9653 ( .A(n13878), .B(n13227), .Z(n12932) );
  CND2X4 U9654 ( .A(n13123), .B(n13128), .Z(n12997) );
  CND2X4 U9655 ( .A(n13123), .B(n15583), .Z(n13124) );
  CND2X4 U9656 ( .A(n12763), .B(n13126), .Z(n12291) );
  CND2X4 U9657 ( .A(n13878), .B(n13128), .Z(n13129) );
  CND2X4 U9658 ( .A(n13100), .B(n12994), .Z(n12175) );
  CND2X4 U9659 ( .A(n13878), .B(n13118), .Z(n12008) );
  CND2X4 U9660 ( .A(n13267), .B(n13126), .Z(n12192) );
  CND2X4 U9661 ( .A(n13267), .B(n13120), .Z(n16425) );
  CND2X4 U9662 ( .A(n13878), .B(n13126), .Z(n16694) );
  CND2X4 U9663 ( .A(n13267), .B(n13877), .Z(n12299) );
  CND2X4 U9664 ( .A(n13100), .B(n13136), .Z(n18028) );
  CND2X4 U9665 ( .A(n13878), .B(n13120), .Z(n12009) );
  CND2X4 U9666 ( .A(n13267), .B(n13128), .Z(n12210) );
  CND2X4 U9667 ( .A(n13878), .B(n12610), .Z(n12202) );
  CND2X4 U9668 ( .A(n13123), .B(n13126), .Z(n12161) );
  CND2X4 U9669 ( .A(n13100), .B(n13877), .Z(n12170) );
  CIVDX1 U9670 ( .A(n12968), .Z0(n12003), .Z1(n17188) );
  CND2X4 U9671 ( .A(n13100), .B(n13120), .Z(n17217) );
  CNIVX4 U9672 ( .A(n11967), .Z(n13493) );
  CND2X4 U9673 ( .A(n13189), .B(n13136), .Z(n13351) );
  CND2X4 U9674 ( .A(n13267), .B(n12610), .Z(n17053) );
  CIVDX1 U9675 ( .A(n12776), .Z0(n12010), .Z1(n12011) );
  CND2X1 U9676 ( .A(n17744), .B(lfsrdin[0]), .Z(n12776) );
  CND2X4 U9677 ( .A(n13267), .B(n13266), .Z(n12012) );
  CIVDX2 U9678 ( .A(n12157), .Z0(n12013), .Z1(n12014) );
  CND2X4 U9679 ( .A(n13100), .B(n12988), .Z(n12401) );
  CIVDX1 U9680 ( .A(n15405), .Z0(n12015), .Z1(n12016) );
  CIVDX1 U9681 ( .A(n12015), .Z0(n13904), .Z1(n15574) );
  CIVDX1 U9682 ( .A(n12015), .Z0(n15403), .Z1(n17031) );
  CIVX8 U9683 ( .A(n17160), .Z(n18017) );
  CIVX2 U9684 ( .A(n12004), .Z(n17423) );
  CND2X2 U9685 ( .A(n17829), .B(lfsrdin[23]), .Z(n12296) );
  CIVDX2 U9686 ( .A(n17721), .Z0(n13994), .Z1(n16179) );
  CNR2X4 U9687 ( .A(n12107), .B(n12102), .Z(n12071) );
  CNIVX1 U9688 ( .A(n12165), .Z(n12572) );
  CND2X4 U9689 ( .A(n18004), .B(n17744), .Z(n12017) );
  CND2X2 U9690 ( .A(n17744), .B(lfsrdin[24]), .Z(n17721) );
  CIVDX4 U9691 ( .A(n12023), .Z0(n12018), .Z1(n12019) );
  CND2X2 U9692 ( .A(n17495), .B(lfsrdin[17]), .Z(n17076) );
  CND2X1 U9693 ( .A(n17959), .B(lfsrdin[16]), .Z(n13449) );
  CIVDX1 U9694 ( .A(n13449), .Z0(n12381), .Z1(n17211) );
  CIVDX2 U9695 ( .A(n14977), .Z0(n14875), .Z1(n12535) );
  CIVDX1 U9696 ( .A(n14977), .Z0(n14868), .Z1(n14645) );
  CIVDX1 U9697 ( .A(n15671), .Z0(n15672) );
  CND2X4 U9698 ( .A(n13123), .B(n12610), .Z(n12598) );
  CIVX2 U9699 ( .A(dataselector[47]), .Z(n14393) );
  CND2X4 U9700 ( .A(n13493), .B(dataselector[25]), .Z(n12214) );
  CNR2IX4 U9701 ( .B(dataselector[21]), .A(n12214), .Z(n12054) );
  CNR2IX2 U9702 ( .B(n14393), .A(n12051), .Z(n12023) );
  CND2X1 U9703 ( .A(n12019), .B(entrophy[8]), .Z(n14998) );
  CND2X4 U9704 ( .A(n12068), .B(dataselector[14]), .Z(n14652) );
  CIVX8 U9705 ( .A(n14652), .Z(n14866) );
  CIVDX2 U9706 ( .A(n12028), .Z0(n12024), .Z1(n12031) );
  CIVX20 U9707 ( .A(rst), .Z(n18257) );
  CND2X4 U9708 ( .A(n16249), .B(n18257), .Z(n14977) );
  CND2X2 U9709 ( .A(n14866), .B(n14875), .Z(n12027) );
  CND2X4 U9710 ( .A(n14033), .B(n14866), .Z(n15335) );
  CIVX2 U9711 ( .A(n15335), .Z(n15274) );
  CAN2X1 U9712 ( .A(dataselector[8]), .B(n18257), .Z(n12025) );
  CND2X2 U9713 ( .A(n12124), .B(n12025), .Z(n15042) );
  CND3XL U9714 ( .A(n15274), .B(n17804), .C(entrophy[11]), .Z(n12026) );
  COAN1X1 U9715 ( .A(n14998), .B(n17763), .C(n12026), .Z(n12063) );
  CIVX2 U9716 ( .A(entrophy[0]), .Z(n17808) );
  CND2X4 U9717 ( .A(n12031), .B(dataselector[21]), .Z(n17805) );
  CIVX2 U9718 ( .A(n14796), .Z(n14392) );
  CND2X2 U9719 ( .A(n17805), .B(n14392), .Z(n12029) );
  CNR2X4 U9720 ( .A(n14782), .B(n12029), .Z(n14454) );
  CND2X2 U9721 ( .A(n15145), .B(n14454), .Z(n14958) );
  CIVX2 U9722 ( .A(dataselector[14]), .Z(n15349) );
  CND2IX4 U9723 ( .B(n14393), .A(n12054), .Z(n13958) );
  CND2X1 U9724 ( .A(n18234), .B(entrophy[29]), .Z(n14894) );
  CIVX2 U9725 ( .A(n14894), .Z(n14879) );
  CND3XL U9726 ( .A(n15043), .B(n17804), .C(n14879), .Z(n12030) );
  COAN1X1 U9727 ( .A(n17808), .B(n14958), .C(n12030), .Z(n12062) );
  CNR2X2 U9728 ( .A(n12214), .B(dataselector[21]), .Z(n12032) );
  CND2X2 U9729 ( .A(n12124), .B(dataselector[47]), .Z(n12043) );
  CNIVX4 U9730 ( .A(n12043), .Z(n14139) );
  CND2X4 U9731 ( .A(n12032), .B(n14139), .Z(n15283) );
  CIVX4 U9732 ( .A(n15283), .Z(n15256) );
  CND2X1 U9733 ( .A(n15256), .B(datain[4]), .Z(n13946) );
  CIVX2 U9734 ( .A(datain[5]), .Z(n14545) );
  CNR2X1 U9735 ( .A(n14796), .B(n14545), .Z(n15160) );
  CIVX1 U9736 ( .A(dataselector[21]), .Z(n14085) );
  CIVX1 U9737 ( .A(n14218), .Z(n12033) );
  CNR2IX2 U9738 ( .B(n14652), .A(n15042), .Z(n15314) );
  CND2X1 U9739 ( .A(n12033), .B(n15314), .Z(n12038) );
  CIVX4 U9740 ( .A(n17805), .Z(n14395) );
  CNIVX4 U9741 ( .A(n12043), .Z(n12034) );
  CIVX8 U9742 ( .A(n12034), .Z(n15302) );
  CND2X2 U9743 ( .A(n14395), .B(n15302), .Z(n14640) );
  CNIVX8 U9744 ( .A(n12214), .Z(n11969) );
  CIVX8 U9745 ( .A(n11969), .Z(n14672) );
  CND2X1 U9746 ( .A(n14672), .B(entrophy[28]), .Z(n15098) );
  CNR2X1 U9747 ( .A(n14640), .B(n15098), .Z(n14956) );
  CIVXL U9748 ( .A(n14956), .Z(n12035) );
  CNR2X4 U9749 ( .A(n17805), .B(dataselector[25]), .Z(n15303) );
  CND2X4 U9750 ( .A(n15303), .B(n15302), .Z(n14969) );
  CIVX4 U9751 ( .A(n14969), .Z(n17759) );
  CND2X1 U9752 ( .A(n17759), .B(entrophy[16]), .Z(n15345) );
  CND4X1 U9753 ( .A(n13946), .B(n12038), .C(n12035), .D(n15345), .Z(n12042) );
  CND2X4 U9754 ( .A(n15302), .B(n17805), .Z(n14633) );
  CNR2X4 U9755 ( .A(n14633), .B(n14782), .Z(n15200) );
  CND2X1 U9756 ( .A(n14084), .B(entrophy[4]), .Z(n14140) );
  CIVX1 U9757 ( .A(n14140), .Z(n12041) );
  CND2X2 U9758 ( .A(n17805), .B(dataselector[47]), .Z(n12036) );
  CNR2X4 U9759 ( .A(n12036), .B(n12214), .Z(n15206) );
  CND2X1 U9760 ( .A(n15206), .B(entrophy[20]), .Z(n12510) );
  CIVX4 U9761 ( .A(n12028), .Z(n12165) );
  CND2XL U9762 ( .A(n17259), .B(scrambler[22]), .Z(n12037) );
  CND2X2 U9763 ( .A(n15303), .B(n14139), .Z(n14132) );
  CND2X1 U9764 ( .A(n14695), .B(datain[5]), .Z(n14827) );
  CND3XL U9765 ( .A(n12510), .B(n12037), .C(n14827), .Z(n12040) );
  COND11X2 U9766 ( .A(n12042), .B(n12041), .C(n12040), .D(n12039), .Z(n12048)
         );
  CNR2X2 U9767 ( .A(n14633), .B(n14782), .Z(n14826) );
  CND2X1 U9768 ( .A(n14826), .B(entrophy[10]), .Z(n14231) );
  CNIVX2 U9769 ( .A(n12043), .Z(n14396) );
  CND2X2 U9770 ( .A(n14395), .B(n14396), .Z(n17809) );
  CND2X2 U9771 ( .A(n17809), .B(n14633), .Z(n14928) );
  CIVX1 U9772 ( .A(n14928), .Z(n14369) );
  CIVX2 U9773 ( .A(entrophy[3]), .Z(n14966) );
  CND2X1 U9774 ( .A(n14695), .B(entrophy[2]), .Z(n15024) );
  CND2X1 U9775 ( .A(n14454), .B(entrophy[31]), .Z(n14909) );
  CND2X1 U9776 ( .A(n14033), .B(entrophy[23]), .Z(n15270) );
  CND2X1 U9777 ( .A(n17759), .B(entrophy[30]), .Z(n14383) );
  CIVX8 U9778 ( .A(n15206), .Z(n15351) );
  COR2XL U9779 ( .A(n15351), .B(n14545), .Z(n12044) );
  CND2X1 U9780 ( .A(n14383), .B(n12044), .Z(n12461) );
  CIVX1 U9781 ( .A(n12461), .Z(n12045) );
  CND2X2 U9782 ( .A(n14875), .B(n14652), .Z(n17785) );
  CANR11X1 U9783 ( .A(n14231), .B(n12046), .C(n12045), .D(n17785), .Z(n12047)
         );
  CNR2IX2 U9784 ( .B(n12048), .A(n12047), .Z(n12061) );
  CND2XL U9785 ( .A(n17804), .B(entrophy[3]), .Z(n15336) );
  CNR2X2 U9786 ( .A(n12266), .B(dataselector[14]), .Z(n12553) );
  CNR2X2 U9787 ( .A(n14788), .B(n14969), .Z(n15306) );
  CND2X4 U9788 ( .A(n17804), .B(dataselector[14]), .Z(n17778) );
  CNR2X2 U9789 ( .A(n14969), .B(n17778), .Z(n17774) );
  CIVX2 U9790 ( .A(n17774), .Z(n15230) );
  CIVX2 U9791 ( .A(entrophy[30]), .Z(n14807) );
  COND2X1 U9792 ( .A(n15336), .B(n14935), .C(n15230), .D(n14807), .Z(n12059)
         );
  CND2X1 U9793 ( .A(n15256), .B(datain[0]), .Z(n14684) );
  CND2X4 U9794 ( .A(n14672), .B(n14396), .Z(n12448) );
  CND2X1 U9795 ( .A(n12214), .B(n15302), .Z(n15299) );
  CND2X2 U9796 ( .A(n12448), .B(n15299), .Z(n14887) );
  CIVX2 U9797 ( .A(entrophy[28]), .Z(n15044) );
  CNR2XL U9798 ( .A(n14395), .B(n15044), .Z(n12049) );
  CND2X1 U9799 ( .A(n12534), .B(n12049), .Z(n12050) );
  CIVX2 U9800 ( .A(n17809), .Z(n17797) );
  CND2X1 U9801 ( .A(n17797), .B(entrophy[0]), .Z(n14781) );
  CNR2X1 U9802 ( .A(n14781), .B(n14672), .Z(n14129) );
  CIVX2 U9803 ( .A(n14129), .Z(n15260) );
  CND2X1 U9804 ( .A(n14857), .B(entrophy[26]), .Z(n14558) );
  CNIVX1 U9805 ( .A(n12051), .Z(n17799) );
  CNR2IX1 U9806 ( .B(datain[0]), .A(n17799), .Z(n14878) );
  CIVX1 U9807 ( .A(n14878), .Z(n12053) );
  CIVX2 U9808 ( .A(entrophy[23]), .Z(n13947) );
  COR2XL U9809 ( .A(n14633), .B(n13947), .Z(n12052) );
  CIVDX2 U9810 ( .A(n12054), .Z0(n12051), .Z1(n15110) );
  CND2X1 U9811 ( .A(n17804), .B(n15349), .Z(n12055) );
  CIVX2 U9812 ( .A(n12055), .Z(n15220) );
  CND2X1 U9813 ( .A(n12057), .B(n12056), .Z(n12058) );
  CNIVX8 U9814 ( .A(n12165), .Z(n17826) );
  CIVX2 U9815 ( .A(n12385), .Z(n12066) );
  CND2X2 U9816 ( .A(n12064), .B(dataselector[1]), .Z(n12596) );
  CNR2IX1 U9817 ( .B(dataselector[31]), .A(n12596), .Z(n12065) );
  CND2X2 U9818 ( .A(n12066), .B(n12065), .Z(n12115) );
  CND2X4 U9819 ( .A(n12092), .B(n16349), .Z(n12112) );
  CND2X2 U9820 ( .A(n12073), .B(dataselector[57]), .Z(n12109) );
  CIVX2 U9821 ( .A(dataselector[31]), .Z(n13479) );
  CIVXL U9822 ( .A(dataselector[53]), .Z(n18244) );
  CNR2X4 U9823 ( .A(n12109), .B(n12074), .Z(n16872) );
  CNR2IX2 U9824 ( .B(dataselector[53]), .A(n16349), .Z(n12069) );
  CIVDX4 U9825 ( .A(n12069), .Z0(n12107) );
  CIVX1 U9826 ( .A(dataselector[1]), .Z(n12070) );
  CNR2IX4 U9827 ( .B(n12070), .A(n12385), .Z(n12085) );
  CND2IX4 U9828 ( .B(n12072), .A(dataselector[31]), .Z(n13780) );
  CIVX2 U9829 ( .A(n13780), .Z(n12091) );
  CIVX8 U9830 ( .A(n16349), .Z(n12080) );
  CND2IX4 U9831 ( .B(dataselector[53]), .A(n12080), .Z(n12101) );
  CNR2X4 U9832 ( .A(n12104), .B(n12101), .Z(n16841) );
  CANR2X1 U9833 ( .A(n12071), .B(Poly4[58]), .C(n16841), .D(Poly12[16]), .Z(
        n12077) );
  CNR2X4 U9834 ( .A(n12115), .B(n12107), .Z(n16865) );
  CIVX2 U9835 ( .A(dataselector[57]), .Z(n18253) );
  CND2X2 U9836 ( .A(n12073), .B(n18253), .Z(n12093) );
  CND2X1 U9837 ( .A(n12091), .B(n12241), .Z(n12096) );
  CNR2X4 U9838 ( .A(n12093), .B(n12096), .Z(n16874) );
  CANR2X1 U9839 ( .A(n16865), .B(poly1_shifted[295]), .C(n16874), .D(
        poly14_shifted[200]), .Z(n12076) );
  CAN2X1 U9840 ( .A(n17755), .B(Poly10[39]), .Z(n16091) );
  CNR2X4 U9841 ( .A(n12093), .B(n12074), .Z(n16862) );
  CNR2X4 U9842 ( .A(n12093), .B(n12108), .Z(n16877) );
  CANR2X1 U9843 ( .A(n16091), .B(n16862), .C(poly9_shifted[67]), .D(n16877), 
        .Z(n12075) );
  CAN4X1 U9844 ( .A(n12078), .B(n12077), .C(n12076), .D(n12075), .Z(n12123) );
  CNR2X2 U9845 ( .A(n12385), .B(n12596), .Z(n12079) );
  CND2X4 U9846 ( .A(n12079), .B(n13479), .Z(n12113) );
  CNR2X4 U9847 ( .A(n12092), .B(n12080), .Z(n12106) );
  CNR2X4 U9848 ( .A(n12113), .B(n12114), .Z(n16855) );
  CIVX2 U9849 ( .A(n12101), .Z(n12082) );
  CAN2X1 U9850 ( .A(n12596), .B(n13780), .Z(n12081) );
  CND2X4 U9851 ( .A(n12385), .B(n12081), .Z(n12105) );
  CNR2IX4 U9852 ( .B(n12082), .A(n12105), .Z(n16837) );
  CANR2X1 U9853 ( .A(n16855), .B(poly14_shifted[118]), .C(poly7_shifted[104]), 
        .D(n16837), .Z(n12090) );
  CNR2X4 U9854 ( .A(n12102), .B(n12112), .Z(n16876) );
  COR2X2 U9855 ( .A(n12113), .B(n12101), .Z(n12083) );
  CIVX8 U9856 ( .A(n12083), .Z(n16839) );
  CANR2X1 U9857 ( .A(n16876), .B(Poly2[41]), .C(n16839), .D(Poly9[22]), .Z(
        n12089) );
  CNR2X4 U9858 ( .A(n12102), .B(n12114), .Z(n16860) );
  CNR2X4 U9859 ( .A(n12104), .B(n12112), .Z(n16843) );
  CANR2X1 U9860 ( .A(n16860), .B(poly1_shifted[160]), .C(n16843), .D(
        poly7_shifted[390]), .Z(n12088) );
  CND2X2 U9861 ( .A(n12085), .B(n13479), .Z(n12110) );
  CNIVX4 U9862 ( .A(n12086), .Z(n16852) );
  CANR2X1 U9863 ( .A(n12084), .B(poly5_shifted[66]), .C(n16852), .D(
        Poly14[194]), .Z(n12087) );
  CAN4X1 U9864 ( .A(n12090), .B(n12089), .C(n12088), .D(n12087), .Z(n12122) );
  CNR2X4 U9865 ( .A(n12112), .B(n12105), .Z(n16840) );
  CND2X1 U9866 ( .A(n12092), .B(n12091), .Z(n12094) );
  CNR2X4 U9867 ( .A(n12093), .B(n12094), .Z(n16838) );
  CANR2X1 U9868 ( .A(n16840), .B(Poly0[156]), .C(n16838), .D(poly9_shifted[60]), .Z(n12100) );
  CNR2X4 U9869 ( .A(n12104), .B(n12114), .Z(n16873) );
  CNR2X4 U9870 ( .A(n12110), .B(n12101), .Z(n16866) );
  CANR2X1 U9871 ( .A(n16873), .B(poly12_shifted[16]), .C(n16866), .D(Poly6[21]), .Z(n12099) );
  CNR2X4 U9872 ( .A(n12107), .B(n12105), .Z(n16850) );
  CNR2X4 U9873 ( .A(n12109), .B(n12094), .Z(n16854) );
  CANR2X1 U9874 ( .A(n16850), .B(poly9_shifted[68]), .C(n16854), .D(Poly5[82]), 
        .Z(n12098) );
  CNR2X1 U9875 ( .A(n12110), .B(n12107), .Z(n12095) );
  CNIVX4 U9876 ( .A(n12095), .Z(n16842) );
  CNR2X4 U9877 ( .A(n12096), .B(n12109), .Z(n16875) );
  CANR2X1 U9878 ( .A(n16842), .B(Poly6[26]), .C(n16875), .D(Poly4[49]), .Z(
        n12097) );
  CAN4X1 U9879 ( .A(n12100), .B(n12099), .C(n12098), .D(n12097), .Z(n12121) );
  CNR2X1 U9880 ( .A(n12102), .B(n12101), .Z(n12103) );
  CNIVX8 U9881 ( .A(n12103), .Z(n16844) );
  CNR2X4 U9882 ( .A(n12104), .B(n12107), .Z(n16867) );
  CANR2X1 U9883 ( .A(n16844), .B(poly5_shifted[45]), .C(n16867), .D(
        poly7_shifted[152]), .Z(n12119) );
  CNR2IX4 U9884 ( .B(n12106), .A(n12105), .Z(n16849) );
  CNR2X4 U9885 ( .A(n12113), .B(n12107), .Z(n16853) );
  CANR2X1 U9886 ( .A(n16849), .B(poly13_shifted[127]), .C(n16853), .D(
        Poly2[67]), .Z(n12118) );
  CNR2X4 U9887 ( .A(n12109), .B(n12108), .Z(n16863) );
  CANR2X1 U9888 ( .A(n16863), .B(poly4_shifted[26]), .C(n16864), .D(
        poly13_shifted[432]), .Z(n12117) );
  CNR2X4 U9889 ( .A(n12113), .B(n12112), .Z(n16861) );
  CNR2X2 U9890 ( .A(n12115), .B(n12114), .Z(n13208) );
  CNIVX4 U9891 ( .A(n13208), .Z(n12872) );
  CANR2X1 U9892 ( .A(n16861), .B(poly7_shifted[102]), .C(n12872), .D(Poly8[67]), .Z(n12116) );
  CAN4X1 U9893 ( .A(n12119), .B(n12118), .C(n12117), .D(n12116), .Z(n12120) );
  CND4X1 U9894 ( .A(n12123), .B(n12122), .C(n12121), .D(n12120), .Z(n12125) );
  CAOR2X1 U9895 ( .A(polydata[13]), .B(n17826), .C(n12125), .D(n16886), .Z(
        n8697) );
  CIVX2 U9896 ( .A(Poly10[32]), .Z(n13731) );
  CNR2X1 U9897 ( .A(n17826), .B(n13731), .Z(n13783) );
  CANR2X1 U9898 ( .A(n16874), .B(poly5_shifted[63]), .C(n16840), .D(n13783), 
        .Z(n12129) );
  CANR2X1 U9899 ( .A(n16865), .B(Poly4[22]), .C(n16860), .D(Poly12[28]), .Z(
        n12128) );
  CANR2X1 U9900 ( .A(n16875), .B(poly9_shifted[48]), .C(n16862), .D(
        poly0_shifted[202]), .Z(n12127) );
  CANR2X1 U9901 ( .A(n16863), .B(Poly10[13]), .C(Poly10[2]), .D(n16837), .Z(
        n12126) );
  CAN4X1 U9902 ( .A(n12129), .B(n12128), .C(n12127), .D(n12126), .Z(n12146) );
  CIVX4 U9903 ( .A(n17160), .Z(n17298) );
  CND2X1 U9904 ( .A(n17298), .B(Poly6[50]), .Z(n13481) );
  CANR2X1 U9905 ( .A(n16838), .B(n13499), .C(poly7_shifted[146]), .D(n12084), 
        .Z(n12133) );
  CANR2X1 U9906 ( .A(n16849), .B(Poly6[15]), .C(n16853), .D(poly11_shifted[15]), .Z(n12132) );
  CANR2X1 U9907 ( .A(n16842), .B(poly11_shifted[29]), .C(n16861), .D(
        poly0_shifted[212]), .Z(n12131) );
  CANR2X1 U9908 ( .A(n16850), .B(poly14_shifted[253]), .C(n16844), .D(
        poly14_shifted[208]), .Z(n12130) );
  CAN4X1 U9909 ( .A(n12133), .B(n12132), .C(n12131), .D(n12130), .Z(n12145) );
  CANR2X1 U9910 ( .A(n16867), .B(poly13_shifted[188]), .C(n16841), .D(
        Poly0[207]), .Z(n12137) );
  CND2X1 U9911 ( .A(n17560), .B(Poly5[112]), .Z(n13417) );
  CIVX2 U9912 ( .A(n13417), .Z(n13586) );
  CANR2X1 U9913 ( .A(n16855), .B(n13586), .C(n12872), .D(poly2_shifted[16]), 
        .Z(n12136) );
  CANR2X1 U9914 ( .A(n12067), .B(poly8_shifted[39]), .C(n16852), .D(Poly2[46]), 
        .Z(n12135) );
  CANR2X1 U9915 ( .A(n16843), .B(poly13_shifted[450]), .C(n16877), .D(Poly8[8]), .Z(n12134) );
  CAN4X1 U9916 ( .A(n12137), .B(n12136), .C(n12135), .D(n12134), .Z(n12144) );
  CANR2X1 U9917 ( .A(n12071), .B(poly0_shifted[215]), .C(n16873), .D(
        Poly11[61]), .Z(n12142) );
  CANR2X1 U9918 ( .A(n16839), .B(Poly6[11]), .C(n16864), .D(poly3_shifted[83]), 
        .Z(n12141) );
  CIVX2 U9919 ( .A(n15648), .Z(n17668) );
  CND2X1 U9920 ( .A(n17668), .B(Poly15[59]), .Z(n16555) );
  CIVXL U9921 ( .A(n16555), .Z(n12138) );
  CANR2X1 U9922 ( .A(n16876), .B(n12138), .C(n16866), .D(poly0_shifted[70]), 
        .Z(n12140) );
  CANR2X1 U9923 ( .A(n16854), .B(Poly10[16]), .C(n16872), .D(
        poly12_shifted[113]), .Z(n12139) );
  CAN4X1 U9924 ( .A(n12142), .B(n12141), .C(n12140), .D(n12139), .Z(n12143) );
  CND4X1 U9925 ( .A(n12146), .B(n12145), .C(n12144), .D(n12143), .Z(n12147) );
  CAOR2X1 U9926 ( .A(polydata[3]), .B(n17259), .C(n12147), .D(n16886), .Z(
        n8687) );
  CENX1 U9927 ( .A(Poly4[51]), .B(n13928), .Z(n15640) );
  CEOX1 U9928 ( .A(Poly4[47]), .B(n15640), .Z(n13140) );
  CEOX2 U9929 ( .A(Poly4[60]), .B(Poly4[56]), .Z(n15651) );
  CENX2 U9930 ( .A(Poly4[55]), .B(Poly4[59]), .Z(n18214) );
  CENX1 U9931 ( .A(Poly4[49]), .B(n18214), .Z(n14613) );
  CENX1 U9932 ( .A(n15651), .B(n14613), .Z(n17326) );
  CENX1 U9933 ( .A(n13140), .B(n17326), .Z(n17219) );
  CIVX1 U9934 ( .A(Poly4[19]), .Z(n12254) );
  CND2XL U9935 ( .A(n17998), .B(n12254), .Z(n12156) );
  CNR2X1 U9936 ( .A(addr[7]), .B(n12158), .Z(n12151) );
  CIVX3 U9937 ( .A(n12191), .Z(n12242) );
  CIVX1 U9938 ( .A(addr[5]), .Z(n12190) );
  CNR2XL U9939 ( .A(addr[4]), .B(n12190), .Z(n12152) );
  CND2X1 U9940 ( .A(n12242), .B(n12152), .Z(n12648) );
  CND2X2 U9941 ( .A(n12648), .B(n17826), .Z(n12250) );
  CIVX2 U9942 ( .A(addr[2]), .Z(n12159) );
  CIVX2 U9943 ( .A(addr[0]), .Z(n12166) );
  CNR2X1 U9944 ( .A(n12166), .B(addr[1]), .Z(n12201) );
  CIVX2 U9945 ( .A(n12201), .Z(n12247) );
  COND1X2 U9946 ( .A(n12277), .B(n12247), .C(n17826), .Z(n13145) );
  CMXI2XL U9947 ( .A0(n12004), .A1(Poly4[36]), .S(n12153), .Z(n12155) );
  CIVX2 U9948 ( .A(n15648), .Z(n17317) );
  CND3XL U9949 ( .A(Poly4[19]), .B(n17317), .C(n17219), .Z(n12154) );
  COND3XL U9950 ( .A(n17219), .B(n12156), .C(n12155), .D(n12154), .Z(n8820) );
  CEOX1 U9951 ( .A(Poly12[58]), .B(Poly12[117]), .Z(n12164) );
  CND2X1 U9952 ( .A(n17668), .B(Poly12[118]), .Z(n14110) );
  CNIVX8 U9953 ( .A(n13493), .Z(n17705) );
  CND2X1 U9954 ( .A(n14107), .B(n12164), .Z(n12163) );
  CND2X1 U9955 ( .A(n17829), .B(lfsrdin[10]), .Z(n12157) );
  CND2IX2 U9956 ( .B(n12158), .A(addr[7]), .Z(n12200) );
  CNR2X2 U9957 ( .A(addr[6]), .B(n12200), .Z(n12183) );
  CND3X1 U9958 ( .A(n12183), .B(addr[5]), .C(addr[4]), .Z(n17967) );
  CND2X2 U9959 ( .A(n17967), .B(n15648), .Z(n13123) );
  CNR2X2 U9960 ( .A(addr[3]), .B(n12159), .Z(n12209) );
  CIVX1 U9961 ( .A(n12209), .Z(n12160) );
  COND1X2 U9962 ( .A(n12404), .B(n12160), .C(n17495), .Z(n13126) );
  CMXI2XL U9963 ( .A0(n12013), .A1(poly12_shifted[90]), .S(n12161), .Z(n12162)
         );
  COND3XL U9964 ( .A(n12164), .B(n14110), .C(n12163), .D(n12162), .Z(n10458)
         );
  CENX1 U9965 ( .A(Poly4[58]), .B(n15640), .Z(n16906) );
  CIVX2 U9966 ( .A(n15673), .Z(n17136) );
  COND1XL U9967 ( .A(n14613), .B(n16906), .C(n17136), .Z(n12168) );
  CNIVX12 U9968 ( .A(n12173), .Z(n17959) );
  COND1X2 U9969 ( .A(n12278), .B(n12277), .C(n17959), .Z(n13136) );
  CND2X4 U9970 ( .A(n12250), .B(n13136), .Z(n18230) );
  CMXI2X1 U9971 ( .A0(n11994), .A1(poly4_shifted[22]), .S(n18230), .Z(n12167)
         );
  COND4CXL U9972 ( .A(n16906), .B(n14613), .C(n12168), .D(n12167), .Z(n8851)
         );
  COND1XL U9973 ( .A(Poly7[401]), .B(Poly7[50]), .C(n18047), .Z(n12172) );
  CNR2X2 U9974 ( .A(addr[4]), .B(addr[5]), .Z(n12268) );
  CND2X1 U9975 ( .A(n12268), .B(n12183), .Z(n12169) );
  CND2X4 U9976 ( .A(n12169), .B(n17495), .Z(n13100) );
  COND1X2 U9977 ( .A(n12356), .B(n12278), .C(n17959), .Z(n13877) );
  CMXI2XL U9978 ( .A0(n18105), .A1(poly7_shifted[74]), .S(n12170), .Z(n12171)
         );
  COND4CXL U9979 ( .A(Poly7[50]), .B(Poly7[401]), .C(n12172), .D(n12171), .Z(
        n10042) );
  CNIVX8 U9980 ( .A(n12173), .Z(n17744) );
  CND2X1 U9981 ( .A(addr[3]), .B(addr[2]), .Z(n12405) );
  CNR2X1 U9982 ( .A(n12405), .B(n12243), .Z(n17964) );
  CIVX2 U9983 ( .A(n17964), .Z(n12174) );
  CND2X2 U9984 ( .A(n17744), .B(n12174), .Z(n12994) );
  CND2X2 U9985 ( .A(n17826), .B(lfsrdin[11]), .Z(n16994) );
  CND2X1 U9986 ( .A(n12175), .B(Poly8[11]), .Z(n12177) );
  CIVX2 U9987 ( .A(n15648), .Z(n16919) );
  CND2X1 U9988 ( .A(n16919), .B(Poly8[93]), .Z(n12176) );
  COND3XL U9989 ( .A(n12175), .B(n16605), .C(n12177), .D(n12176), .Z(n11390)
         );
  COND1XL U9990 ( .A(Poly7[408]), .B(Poly7[242]), .C(n17998), .Z(n12179) );
  CND2X4 U9991 ( .A(n13100), .B(n13126), .Z(n17574) );
  CMXI2XL U9992 ( .A0(n18105), .A1(poly7_shifted[266]), .S(n17574), .Z(n12178)
         );
  COND4CXL U9993 ( .A(Poly7[242]), .B(Poly7[408]), .C(n12179), .D(n12178), .Z(
        n9850) );
  CND2X1 U9994 ( .A(n12005), .B(n17829), .Z(n18131) );
  COND1X2 U9995 ( .A(n12356), .B(n12243), .C(n17826), .Z(n13118) );
  CND2X2 U9996 ( .A(n12250), .B(n13118), .Z(n17589) );
  COND1XL U9997 ( .A(Poly5[80]), .B(Poly5[115]), .C(n17288), .Z(n12181) );
  CND3X1 U9998 ( .A(n12242), .B(addr[4]), .C(addr[5]), .Z(n18019) );
  CND2X2 U9999 ( .A(n18019), .B(n17160), .Z(n12704) );
  CMXI2XL U10000 ( .A0(n18105), .A1(Poly5[94]), .S(n17942), .Z(n12180) );
  COND4CXL U10001 ( .A(Poly5[115]), .B(Poly5[80]), .C(n12181), .D(n12180), .Z(
        n11432) );
  CIVXL U10002 ( .A(addr[4]), .Z(n12182) );
  CND2XL U10003 ( .A(addr[5]), .B(n12182), .Z(n12184) );
  CIVX2 U10004 ( .A(n12183), .Z(n12260) );
  COND1X2 U10005 ( .A(n12184), .B(n12260), .C(n17959), .Z(n12396) );
  COND1X2 U10006 ( .A(n12404), .B(n12277), .C(n17959), .Z(n13093) );
  CND2X1 U10007 ( .A(n12185), .B(poly11_shifted[19]), .Z(n12186) );
  CENX1 U10008 ( .A(Poly11[83]), .B(Poly11[75]), .Z(n17628) );
  COND3XL U10009 ( .A(n12185), .B(n12005), .C(n12186), .D(n15246), .Z(n11185)
         );
  COND1XL U10010 ( .A(Poly5[116]), .B(Poly5[81]), .C(n17238), .Z(n12188) );
  CMXI2XL U10011 ( .A0(n14436), .A1(Poly5[95]), .S(n17942), .Z(n12187) );
  COND4CXL U10012 ( .A(Poly5[81]), .B(Poly5[116]), .C(n12188), .D(n12187), .Z(
        n11431) );
  CND2X2 U10013 ( .A(n17829), .B(lfsrdin[14]), .Z(n12764) );
  CND2X1 U10014 ( .A(n18017), .B(Poly3[71]), .Z(n13766) );
  CIVX1 U10015 ( .A(Poly3[71]), .Z(n12652) );
  CND2X1 U10016 ( .A(n17317), .B(n12652), .Z(n12614) );
  CMX2GX1 U10017 ( .GN(n18160), .A0(n13766), .A1(n12614), .S(Poly3[32]), .Z(
        n12189) );
  CIVX2 U10018 ( .A(Poly3[46]), .Z(n12615) );
  CMXI2X1 U10019 ( .A0(n12189), .A1(n12615), .S(n17262), .Z(n8894) );
  COND1XL U10020 ( .A(Poly1[343]), .B(Poly1[232]), .C(n16488), .Z(n12194) );
  CND2X2 U10021 ( .A(addr[4]), .B(n12190), .Z(n12261) );
  CMXI2XL U10022 ( .A0(n18176), .A1(poly1_shifted[254]), .S(n12192), .Z(n12193) );
  COND4CXL U10023 ( .A(Poly1[232]), .B(Poly1[343]), .C(n12194), .D(n12193), 
        .Z(n9114) );
  COND1XL U10024 ( .A(Poly12[112]), .B(Poly12[82]), .C(n18234), .Z(n12196) );
  CAN2X4 U10025 ( .A(n13123), .B(n13227), .Z(n18001) );
  CMXI2XL U10026 ( .A0(poly12_shifted[114]), .A1(n12415), .S(n18001), .Z(
        n12195) );
  COND4CXL U10027 ( .A(Poly12[82]), .B(Poly12[112]), .C(n12196), .D(n12195), 
        .Z(n10434) );
  CIVX2 U10028 ( .A(n15648), .Z(n17063) );
  COND1XL U10029 ( .A(Poly12[117]), .B(Poly12[87]), .C(n17063), .Z(n12198) );
  CMXI2XL U10030 ( .A0(poly12_shifted[119]), .A1(n18138), .S(n18001), .Z(
        n12197) );
  COND4CXL U10031 ( .A(Poly12[87]), .B(Poly12[117]), .C(n12198), .D(n12197), 
        .Z(n10429) );
  CIVXL U10032 ( .A(Poly12[123]), .Z(n12199) );
  CND2X1 U10033 ( .A(n17744), .B(lfsrdin[13]), .Z(n12949) );
  CIVX2 U10034 ( .A(n12949), .Z(n18219) );
  CEOXL U10035 ( .A(Poly14[298]), .B(Poly14[206]), .Z(n12205) );
  COND1XL U10036 ( .A(Poly14[292]), .B(n12205), .C(n17099), .Z(n12204) );
  CND2X1 U10037 ( .A(n12201), .B(n12209), .Z(n12953) );
  CND2X2 U10038 ( .A(n12953), .B(n17744), .Z(n12610) );
  CMXI2XL U10039 ( .A0(n18105), .A1(poly14_shifted[238]), .S(n12202), .Z(
        n12203) );
  COND4CXL U10040 ( .A(n12205), .B(Poly14[292]), .C(n12204), .D(n12203), .Z(
        n10183) );
  CIVX1 U10041 ( .A(poly7_shifted[361]), .Z(n14609) );
  COND1XL U10042 ( .A(n17259), .B(n14609), .C(n12002), .Z(n12207) );
  CMX2XL U10043 ( .A0(n12207), .A1(poly7_shifted[373]), .S(n12206), .Z(n9743)
         );
  CNR2X1 U10044 ( .A(n14361), .B(n13783), .Z(n12208) );
  CIVX2 U10045 ( .A(Poly10[1]), .Z(n16094) );
  COND1X4 U10046 ( .A(n12356), .B(n12247), .C(n17959), .Z(n13266) );
  CIVX4 U10047 ( .A(n13782), .Z(n17962) );
  CMXI2XL U10048 ( .A0(n12208), .A1(n16094), .S(n17962), .Z(n11102) );
  CND2X1 U10049 ( .A(n18234), .B(Poly10[33]), .Z(n13756) );
  CND2X1 U10050 ( .A(n17751), .B(n17744), .Z(n18185) );
  CND2X2 U10051 ( .A(n12649), .B(n17826), .Z(n13128) );
  CNR2X1 U10052 ( .A(n18048), .B(n16700), .Z(n13660) );
  CIVX2 U10053 ( .A(n13660), .Z(n18193) );
  COND1X2 U10054 ( .A(n12243), .B(n12277), .C(n17744), .Z(n12988) );
  CND2X1 U10055 ( .A(n17959), .B(lfsrdin[15]), .Z(n16248) );
  CNIVX8 U10056 ( .A(n16248), .Z(n17196) );
  CND2X1 U10057 ( .A(n17196), .B(n17959), .Z(n18163) );
  COND1XL U10058 ( .A(poly15_shifted[15]), .B(n18206), .C(n18163), .Z(n12213)
         );
  CIVX2 U10059 ( .A(Poly15[15]), .Z(n13419) );
  COND1X1 U10060 ( .A(n12405), .B(n12247), .C(n17495), .Z(n12991) );
  CND2X1 U10061 ( .A(n13878), .B(n12991), .Z(n12212) );
  CMXI2X1 U10062 ( .A0(n12213), .A1(n13419), .S(n18044), .Z(n9622) );
  CND2X1 U10063 ( .A(n17607), .B(datain[6]), .Z(n14644) );
  CIVXL U10064 ( .A(n14644), .Z(n12215) );
  CAN2X1 U10065 ( .A(n15206), .B(n15349), .Z(n14976) );
  CIVDX2 U10066 ( .A(n12214), .Z0(n14782), .Z1(n14687) );
  CND2X1 U10067 ( .A(n14928), .B(n14687), .Z(n14451) );
  COND3XL U10068 ( .A(n12215), .B(n14976), .C(n14451), .D(n15314), .Z(n12220)
         );
  CNR2X2 U10069 ( .A(n14640), .B(dataselector[14]), .Z(n15101) );
  CANR4CX1 U10070 ( .A(entrophy[4]), .B(n15101), .C(n15302), .D(n11969), .Z(
        n12219) );
  CANR2X1 U10071 ( .A(n11971), .B(datain[0]), .C(entrophy[5]), .D(n17787), .Z(
        n12218) );
  CNR2X4 U10072 ( .A(n17778), .B(n12520), .Z(n17812) );
  CIVX2 U10073 ( .A(entrophy[14]), .Z(n14871) );
  CNR2X1 U10074 ( .A(n15283), .B(n14871), .Z(n14134) );
  CND2X2 U10075 ( .A(n14875), .B(n12553), .Z(n15293) );
  CND2X1 U10076 ( .A(n15293), .B(n17778), .Z(n14693) );
  CANR2X1 U10077 ( .A(n17812), .B(entrophy[16]), .C(n14134), .D(n14693), .Z(
        n12217) );
  COND3X1 U10078 ( .A(n12220), .B(n12219), .C(n12218), .D(n12217), .Z(n12221)
         );
  CIVX2 U10079 ( .A(n12221), .Z(n12240) );
  CND2X1 U10080 ( .A(n14652), .B(n14393), .Z(n12456) );
  CNR3X2 U10081 ( .A(n11969), .B(n12456), .C(n17805), .Z(n15354) );
  CIVX2 U10082 ( .A(entrophy[20]), .Z(n14387) );
  CANR2X1 U10083 ( .A(n15354), .B(entrophy[12]), .C(n14864), .D(n13945), .Z(
        n12552) );
  CNR2X1 U10084 ( .A(n12552), .B(n15334), .Z(n12232) );
  CND2X1 U10085 ( .A(n15319), .B(entrophy[28]), .Z(n15252) );
  CIVX2 U10086 ( .A(n15351), .Z(n14540) );
  CND2X1 U10087 ( .A(n14540), .B(entrophy[7]), .Z(n14845) );
  CIVX2 U10088 ( .A(entrophy[5]), .Z(n14886) );
  CNR2X1 U10089 ( .A(n12018), .B(n14886), .Z(n15286) );
  CND2X1 U10090 ( .A(n14680), .B(datain[4]), .Z(n15329) );
  CND2XL U10091 ( .A(n17759), .B(entrophy[17]), .Z(n12222) );
  CND2X1 U10092 ( .A(n14695), .B(entrophy[24]), .Z(n15097) );
  CND2X1 U10093 ( .A(n14826), .B(entrophy[29]), .Z(n15114) );
  CIVX1 U10094 ( .A(n15114), .Z(n12228) );
  CND2X1 U10095 ( .A(n14695), .B(datain[1]), .Z(n14075) );
  CIVX2 U10096 ( .A(datain[7]), .Z(n15339) );
  CNR2X1 U10097 ( .A(n14472), .B(n15339), .Z(n14631) );
  CNR2IX1 U10098 ( .B(n14075), .A(n14631), .Z(n12226) );
  CND2X1 U10099 ( .A(n14540), .B(entrophy[22]), .Z(n17793) );
  CND2X2 U10100 ( .A(n17759), .B(entrophy[13]), .Z(n15208) );
  CND2X1 U10101 ( .A(n14454), .B(datain[3]), .Z(n14415) );
  CND2X1 U10102 ( .A(n15208), .B(n14415), .Z(n12515) );
  CIVX1 U10103 ( .A(n12515), .Z(n12225) );
  CND2X1 U10104 ( .A(n12019), .B(entrophy[31]), .Z(n12224) );
  CND4X1 U10105 ( .A(n12226), .B(n17793), .C(n12225), .D(n12224), .Z(n12227)
         );
  CIVX2 U10106 ( .A(n15293), .Z(n15346) );
  COND1X1 U10107 ( .A(n12228), .B(n12227), .C(n15346), .Z(n12229) );
  COND1X1 U10108 ( .A(n12230), .B(n17763), .C(n12229), .Z(n12231) );
  CNR2X2 U10109 ( .A(n12232), .B(n12231), .Z(n12239) );
  CNR2X1 U10110 ( .A(n15283), .B(n15339), .Z(n14697) );
  CND2XL U10111 ( .A(n14697), .B(n14652), .Z(n14421) );
  CIVX2 U10112 ( .A(entrophy[21]), .Z(n14561) );
  CNR2X1 U10113 ( .A(n14226), .B(n14561), .Z(n14588) );
  CIVDX3 U10114 ( .A(n12018), .Z0(n14033), .Z1(n14546) );
  CIVX2 U10115 ( .A(entrophy[6]), .Z(n14908) );
  CNR2X1 U10116 ( .A(n14546), .B(n14908), .Z(n14985) );
  CIVX2 U10117 ( .A(datain[2]), .Z(n14659) );
  CNR2X1 U10118 ( .A(n13958), .B(n14659), .Z(n15295) );
  COND11X1 U10119 ( .A(n14588), .B(n14985), .C(n15295), .D(n12216), .Z(n12236)
         );
  CIVX2 U10120 ( .A(entrophy[15]), .Z(n17784) );
  CIVX2 U10121 ( .A(n15314), .Z(n15170) );
  CND2XL U10122 ( .A(n17744), .B(scrambler[21]), .Z(n12233) );
  COND11X1 U10123 ( .A(n17784), .B(n15170), .C(n14226), .D(n12233), .Z(n12234)
         );
  CANR1XL U10124 ( .A(entrophy[17]), .B(n17774), .C(n12234), .Z(n12235) );
  COND3X1 U10125 ( .A(n14421), .B(n15334), .C(n12236), .D(n12235), .Z(n12237)
         );
  CIVX2 U10126 ( .A(n12237), .Z(n12238) );
  CND3XL U10127 ( .A(n12240), .B(n12239), .C(n12238), .Z(n8721) );
  CENX1 U10128 ( .A(dataselector[59]), .B(dataselector[58]), .Z(n16384) );
  CIVX1 U10129 ( .A(n16384), .Z(n18245) );
  COND1XL U10130 ( .A(n18245), .B(n12241), .C(n11978), .Z(n12244) );
  CND2X4 U10131 ( .A(n12242), .B(n12268), .Z(n18184) );
  CNR3X2 U10132 ( .A(n12243), .B(n12356), .C(n18184), .Z(n12364) );
  CNR2X1 U10133 ( .A(n12364), .B(n18017), .Z(n13882) );
  CIVX4 U10134 ( .A(n18252), .Z(n16350) );
  CMXI2X1 U10135 ( .A0(n12244), .A1(dataselector[60]), .S(n16350), .Z(n12245)
         );
  COND11XL U10136 ( .A(dataselector[53]), .B(n17826), .C(n16384), .D(n12245), 
        .Z(n8735) );
  CENX1 U10137 ( .A(Poly0[161]), .B(Poly0[213]), .Z(n12246) );
  COND1XL U10138 ( .A(n12246), .B(n17959), .C(n17661), .Z(n12249) );
  COR2X1 U10139 ( .A(n12277), .B(n12247), .Z(n12248) );
  CNR2X4 U10140 ( .A(n18184), .B(n12248), .Z(n15960) );
  CMX2XL U10141 ( .A0(n12249), .A1(poly0_shifted[197]), .S(n15671), .Z(n9398)
         );
  CND2XL U10142 ( .A(n13493), .B(Poly3[79]), .Z(n13371) );
  CND2X1 U10143 ( .A(n15737), .B(poly3_shifted[23]), .Z(n12251) );
  COND4CX1 U10144 ( .A(n12002), .B(n13371), .C(n15737), .D(n12251), .Z(n8931)
         );
  CND2X1 U10145 ( .A(n12396), .B(n12988), .Z(n13421) );
  CIVX4 U10146 ( .A(n11998), .Z(n17683) );
  CND2X1 U10147 ( .A(n17683), .B(Poly11[38]), .Z(n12253) );
  CENX1 U10148 ( .A(Poly11[85]), .B(Poly11[77]), .Z(n15385) );
  CNR2X1 U10149 ( .A(n17744), .B(n15385), .Z(n16415) );
  CIVX1 U10150 ( .A(n15385), .Z(n14014) );
  CNR2X1 U10151 ( .A(n17744), .B(n14014), .Z(n13488) );
  CMXI2XL U10152 ( .A0(n16415), .A1(n13488), .S(Poly11[23]), .Z(n12252) );
  COND3XL U10153 ( .A(n17683), .B(n17757), .C(n12253), .D(n12252), .Z(n11151)
         );
  CND2X1 U10154 ( .A(n17673), .B(n17259), .Z(n18175) );
  COND1XL U10155 ( .A(poly4_shifted[19]), .B(n18176), .C(n18175), .Z(n12255)
         );
  CMXI2XL U10156 ( .A0(n12255), .A1(n12254), .S(n18230), .Z(n8837) );
  CIVX8 U10157 ( .A(n15648), .Z(n17538) );
  CENX1 U10158 ( .A(Poly2[68]), .B(Poly2[61]), .Z(n12256) );
  CIVX2 U10159 ( .A(n17310), .Z(n17313) );
  CIVX8 U10160 ( .A(n15673), .Z(n17535) );
  CND2X1 U10161 ( .A(n17535), .B(n12256), .Z(n17307) );
  CIVX2 U10162 ( .A(n17307), .Z(n13647) );
  CMXI2X1 U10163 ( .A0(n17313), .A1(n13647), .S(Poly2[49]), .Z(n12258) );
  COND1X1 U10164 ( .A(n12405), .B(n12278), .C(n15648), .Z(n12395) );
  CMXI2XL U10165 ( .A0(n18228), .A1(Poly2[61]), .S(n17306), .Z(n12257) );
  CND2XL U10166 ( .A(n12258), .B(n12257), .Z(n8949) );
  CND2X1 U10167 ( .A(n17959), .B(lfsrdin[21]), .Z(n12273) );
  CND2X1 U10168 ( .A(n17036), .B(n17826), .Z(n18085) );
  CND2X1 U10169 ( .A(n12185), .B(poly11_shifted[26]), .Z(n12259) );
  CND2X1 U10170 ( .A(n17755), .B(Poly11[82]), .Z(n13507) );
  COND3XL U10171 ( .A(n12185), .B(n16605), .C(n12259), .D(n13507), .Z(n11178)
         );
  CND2X2 U10172 ( .A(n17959), .B(lfsrdin[25]), .Z(n17123) );
  COR2XL U10173 ( .A(Poly12[124]), .B(Poly12[94]), .Z(n12263) );
  CND2XL U10174 ( .A(n17453), .B(n12263), .Z(n12265) );
  CMXI2XL U10175 ( .A0(poly12_shifted[126]), .A1(n18160), .S(n18001), .Z(
        n12264) );
  COND4CX1 U10176 ( .A(Poly12[94]), .B(Poly12[124]), .C(n12265), .D(n12264), 
        .Z(n10422) );
  CND2X1 U10177 ( .A(n17714), .B(Poly15[49]), .Z(n14525) );
  CND2X1 U10178 ( .A(n18044), .B(poly15_shifted[19]), .Z(n12267) );
  COND4CXL U10179 ( .A(n12005), .B(n14525), .C(n18044), .D(n12267), .Z(n9633)
         );
  CND2X1 U10180 ( .A(n17718), .B(n17744), .Z(n18137) );
  CND2IX1 U10181 ( .B(n12269), .A(n12268), .Z(n18004) );
  CND2X1 U10182 ( .A(n12017), .B(n12395), .Z(n12270) );
  CANR2X1 U10183 ( .A(n17990), .B(poly13_shifted[473]), .C(n18234), .D(
        poly13_shifted[459]), .Z(n12271) );
  COND1XL U10184 ( .A(n16605), .B(n17990), .C(n12271), .Z(n10601) );
  CANR2X1 U10185 ( .A(n17990), .B(poly13_shifted[468]), .C(n17449), .D(
        poly13_shifted[454]), .Z(n12272) );
  COND1XL U10186 ( .A(n16779), .B(n17990), .C(n12272), .Z(n10606) );
  CND2X1 U10187 ( .A(n12704), .B(n13877), .Z(n17928) );
  CIVDX2 U10188 ( .A(n17928), .Z0(n15613), .Z1(n17930) );
  CND2XL U10189 ( .A(n17930), .B(poly5_shifted[35]), .Z(n12275) );
  CND2XL U10190 ( .A(n17545), .B(poly5_shifted[21]), .Z(n12274) );
  COND3XL U10191 ( .A(n17932), .B(n12006), .C(n12275), .D(n12274), .Z(n11505)
         );
  CENX1 U10192 ( .A(Poly0[117]), .B(Poly0[216]), .Z(n12276) );
  COND1XL U10193 ( .A(n12276), .B(n17959), .C(n16939), .Z(n12280) );
  CIVX2 U10194 ( .A(n17160), .Z(n17607) );
  CNR3X1 U10195 ( .A(n12278), .B(n12277), .C(n18184), .Z(n12279) );
  CNR2X4 U10196 ( .A(n17607), .B(n14441), .Z(n17671) );
  CMX2XL U10197 ( .A0(n12280), .A1(poly0_shifted[153]), .S(n17671), .Z(n9442)
         );
  CND2X2 U10198 ( .A(n18184), .B(n17744), .Z(n12763) );
  CND2X4 U10199 ( .A(n12763), .B(n12994), .Z(n18180) );
  CND2X1 U10200 ( .A(n13418), .B(n17959), .Z(n18104) );
  CND2X1 U10201 ( .A(n17721), .B(n17495), .Z(n18091) );
  CIVX8 U10202 ( .A(n18228), .Z(n17185) );
  CND2X1 U10203 ( .A(n17185), .B(n17959), .Z(n18227) );
  CND2X1 U10204 ( .A(n11978), .B(n17959), .Z(n18224) );
  CND2X1 U10205 ( .A(n17305), .B(n17959), .Z(n18094) );
  CND2X1 U10206 ( .A(n17741), .B(n15673), .Z(n18098) );
  CND2X1 U10207 ( .A(n17753), .B(n17744), .Z(n18088) );
  CIVX1 U10208 ( .A(Poly12[119]), .Z(n18000) );
  CAN2X1 U10209 ( .A(n17620), .B(n18000), .Z(n17995) );
  COND1XL U10210 ( .A(Poly2[30]), .B(Poly2[66]), .C(n17178), .Z(n12282) );
  CMXI2XL U10211 ( .A0(n12013), .A1(Poly2[42]), .S(n17306), .Z(n12281) );
  COND4CXL U10212 ( .A(Poly2[66]), .B(Poly2[30]), .C(n12282), .D(n12281), .Z(
        n8968) );
  CIVX2 U10213 ( .A(n12001), .Z(n17208) );
  CND2XL U10214 ( .A(n17942), .B(poly5_shifted[87]), .Z(n12284) );
  CND2XL U10215 ( .A(n17266), .B(poly5_shifted[73]), .Z(n12283) );
  COND3XL U10216 ( .A(n17942), .B(n17208), .C(n12284), .D(n12283), .Z(n11453)
         );
  CND2X1 U10217 ( .A(n17757), .B(n17495), .Z(n18117) );
  CIVXL U10218 ( .A(poly8_shifted[38]), .Z(n12285) );
  CND2IX1 U10219 ( .B(n14754), .A(n12285), .Z(n12286) );
  CND2X1 U10220 ( .A(n18117), .B(n12286), .Z(n12289) );
  CND2X1 U10221 ( .A(n12287), .B(poly8_shifted[52]), .Z(n12288) );
  COND1XL U10222 ( .A(n12289), .B(n12287), .C(n12288), .Z(n11363) );
  CND2X2 U10223 ( .A(n17495), .B(lfsrdin[20]), .Z(n16391) );
  CND2X1 U10224 ( .A(n16391), .B(n17744), .Z(n18200) );
  COND1XL U10225 ( .A(poly1_shifted[20]), .B(n18082), .C(n18200), .Z(n12290)
         );
  CIVX2 U10226 ( .A(Poly1[20]), .Z(n18179) );
  CMXI2XL U10227 ( .A0(n12290), .A1(n18179), .S(n18180), .Z(n9337) );
  CIVX2 U10228 ( .A(n17259), .Z(n17156) );
  COND1XL U10229 ( .A(Poly2[68]), .B(Poly2[41]), .C(n17156), .Z(n12293) );
  CMXI2X1 U10230 ( .A0(n18241), .A1(Poly2[53]), .S(n17306), .Z(n12292) );
  COND4CX1 U10231 ( .A(Poly2[41]), .B(Poly2[68]), .C(n12293), .D(n12292), .Z(
        n8957) );
  COND1XL U10232 ( .A(Poly2[67]), .B(Poly2[40]), .C(n16919), .Z(n12295) );
  CMXI2XL U10233 ( .A0(n18082), .A1(Poly2[52]), .S(n17306), .Z(n12294) );
  COND4CXL U10234 ( .A(Poly2[40]), .B(Poly2[67]), .C(n12295), .D(n12294), .Z(
        n8958) );
  CIVX1 U10235 ( .A(poly0_shifted[87]), .Z(n13679) );
  COND1XL U10236 ( .A(n17744), .B(n13679), .C(n12000), .Z(n12297) );
  CMX2XL U10237 ( .A0(n12297), .A1(poly0_shifted[105]), .S(n12291), .Z(n9490)
         );
  CND2X1 U10238 ( .A(n12296), .B(n17826), .Z(n18203) );
  CIVDXL U10239 ( .A(n17123), .Z0(n17934), .Z1(n11997) );
  COND1XL U10240 ( .A(poly1_shifted[25]), .B(n17934), .C(n18196), .Z(n12298)
         );
  CIVX1 U10241 ( .A(Poly1[25]), .Z(n13717) );
  CMXI2XL U10242 ( .A0(n12298), .A1(n13717), .S(n18180), .Z(n9332) );
  CND2X1 U10243 ( .A(n16947), .B(Poly1[339]), .Z(n13223) );
  COAN1XL U10244 ( .A(Poly1[23]), .B(n13223), .C(n16303), .Z(n12301) );
  CANR2X1 U10245 ( .A(n12299), .B(poly1_shifted[45]), .C(Poly1[23]), .D(n13362), .Z(n12300) );
  COND1XL U10246 ( .A(n12301), .B(n12299), .C(n12300), .Z(n9323) );
  COND1XL U10247 ( .A(Poly7[401]), .B(Poly7[235]), .C(n18047), .Z(n12303) );
  CMXI2XL U10248 ( .A0(n11999), .A1(poly7_shifted[259]), .S(n17574), .Z(n12302) );
  COND4CXL U10249 ( .A(Poly7[235]), .B(Poly7[401]), .C(n12303), .D(n12302), 
        .Z(n9857) );
  CND2X1 U10250 ( .A(n13267), .B(n13136), .Z(n12304) );
  CNIVX8 U10251 ( .A(n12304), .Z(n18198) );
  CANR2XL U10252 ( .A(n18198), .B(poly1_shifted[310]), .C(poly1_shifted[299]), 
        .D(n18017), .Z(n12305) );
  COND1XL U10253 ( .A(n16605), .B(n18198), .C(n12305), .Z(n9058) );
  CND2X4 U10254 ( .A(n13267), .B(n13227), .Z(n18191) );
  CANR2X1 U10255 ( .A(n18191), .B(poly1_shifted[267]), .C(n17613), .D(
        poly1_shifted[256]), .Z(n12306) );
  COND1XL U10256 ( .A(n12011), .B(n18191), .C(n12306), .Z(n9101) );
  CANR2X1 U10257 ( .A(n17332), .B(poly1_shifted[342]), .C(n17552), .D(
        poly1_shifted[331]), .Z(n12307) );
  COND1XL U10258 ( .A(n16605), .B(n17332), .C(n12307), .Z(n9026) );
  CANR2X1 U10259 ( .A(n12192), .B(poly1_shifted[263]), .C(n17094), .D(
        poly1_shifted[252]), .Z(n12308) );
  COND1XL U10260 ( .A(n11978), .B(n12192), .C(n12308), .Z(n9105) );
  CANR2X1 U10261 ( .A(n17053), .B(Poly1[201]), .C(n17238), .D(
        poly1_shifted[201]), .Z(n12309) );
  COND1XL U10262 ( .A(n17208), .B(n17053), .C(n12309), .Z(n9156) );
  CIVX2 U10263 ( .A(n17160), .Z(n16947) );
  CND2X1 U10264 ( .A(n16947), .B(Poly15[48]), .Z(n13420) );
  CND2X1 U10265 ( .A(n18044), .B(poly15_shifted[18]), .Z(n12310) );
  COND4CXL U10266 ( .A(n13275), .B(n13420), .C(n18044), .D(n12310), .Z(n9634)
         );
  CND2X1 U10267 ( .A(n18044), .B(Poly15[14]), .Z(n12311) );
  COND4CXL U10268 ( .A(n16555), .B(n17699), .C(n18044), .D(n12311), .Z(n9623)
         );
  CIVX2 U10269 ( .A(n15648), .Z(n16700) );
  CND2X1 U10270 ( .A(n16700), .B(Poly15[54]), .Z(n16740) );
  CND2X1 U10271 ( .A(n18044), .B(poly15_shifted[24]), .Z(n12312) );
  COND4CXL U10272 ( .A(n16740), .B(n12002), .C(n18044), .D(n12312), .Z(n9628)
         );
  CND2X1 U10273 ( .A(n12211), .B(poly2_shifted[15]), .Z(n12313) );
  COND3XL U10274 ( .A(n12211), .B(n13275), .C(n12313), .D(n17310), .Z(n9007)
         );
  CANR2X1 U10275 ( .A(n16861), .B(Poly12[27]), .C(n16875), .D(Poly10[10]), .Z(
        n12317) );
  CANR2X1 U10276 ( .A(n16842), .B(poly5_shifted[58]), .C(n16865), .D(
        poly9_shifted[59]), .Z(n12316) );
  CANR2X1 U10277 ( .A(n12067), .B(poly13_shifted[154]), .C(poly14_shifted[178]), .D(n16849), .Z(n12315) );
  CANR2X1 U10278 ( .A(n16840), .B(poly5_shifted[26]), .C(poly10_shifted[18]), 
        .D(n12872), .Z(n12314) );
  CAN4X1 U10279 ( .A(n12317), .B(n12316), .C(n12315), .D(n12314), .Z(n12333)
         );
  CANR2X1 U10280 ( .A(n16874), .B(Poly8[2]), .C(poly13_shifted[81]), .D(n16837), .Z(n12321) );
  CANR2X1 U10281 ( .A(n16854), .B(Poly11[78]), .C(n16843), .D(Poly11[35]), .Z(
        n12320) );
  CANR2X1 U10282 ( .A(n16844), .B(Poly10[15]), .C(n16876), .D(Poly6[12]), .Z(
        n12319) );
  CANR2X1 U10283 ( .A(n12071), .B(poly3_shifted[44]), .C(n16860), .D(
        poly14_shifted[171]), .Z(n12318) );
  CAN4X1 U10284 ( .A(n12321), .B(n12320), .C(n12319), .D(n12318), .Z(n12332)
         );
  CANR2X1 U10285 ( .A(n16863), .B(poly0_shifted[196]), .C(n12084), .D(
        poly14_shifted[77]), .Z(n12325) );
  CANR2X1 U10286 ( .A(n16872), .B(Poly7[178]), .C(n16877), .D(
        poly5_shifted[82]), .Z(n12324) );
  CANR2X1 U10287 ( .A(n16855), .B(Poly2[24]), .C(n16866), .D(Poly4[25]), .Z(
        n12323) );
  CANR2X1 U10288 ( .A(n16838), .B(poly14_shifted[234]), .C(n16841), .D(
        Poly6[20]), .Z(n12322) );
  CAN4X1 U10289 ( .A(n12325), .B(n12324), .C(n12323), .D(n12322), .Z(n12331)
         );
  CANR2X1 U10290 ( .A(n16850), .B(poly1_shifted[256]), .C(poly3_shifted[79]), 
        .D(n16867), .Z(n12329) );
  CANR2X1 U10291 ( .A(n16864), .B(Poly12[95]), .C(n16862), .D(Poly15[14]), .Z(
        n12328) );
  CANR2X1 U10292 ( .A(n16839), .B(Poly5[114]), .C(n16852), .D(
        poly0_shifted[87]), .Z(n12327) );
  CANR2X1 U10293 ( .A(n16873), .B(poly8_shifted[47]), .C(n16853), .D(
        poly8_shifted[36]), .Z(n12326) );
  CAN4X1 U10294 ( .A(n12329), .B(n12328), .C(n12327), .D(n12326), .Z(n12330)
         );
  CND4X1 U10295 ( .A(n12333), .B(n12332), .C(n12331), .D(n12330), .Z(n12334)
         );
  CAOR2X1 U10296 ( .A(polydata[12]), .B(n17744), .C(n12334), .D(n16886), .Z(
        n8696) );
  CANR2X1 U10297 ( .A(n16860), .B(poly7_shifted[58]), .C(n16866), .D(
        Poly12[64]), .Z(n12338) );
  CND2X1 U10298 ( .A(n17607), .B(Poly15[58]), .Z(n14515) );
  CIVX1 U10299 ( .A(n14515), .Z(n13036) );
  CANR2X1 U10300 ( .A(n16852), .B(n13036), .C(n16843), .D(poly4_shifted[25]), 
        .Z(n12337) );
  CANR2X1 U10301 ( .A(n16850), .B(poly12_shifted[20]), .C(n16876), .D(
        poly0_shifted[164]), .Z(n12336) );
  CANR2X1 U10302 ( .A(n16874), .B(poly1_shifted[305]), .C(Poly11[71]), .D(
        n16837), .Z(n12335) );
  CAN4X1 U10303 ( .A(n12338), .B(n12337), .C(n12336), .D(n12335), .Z(n12354)
         );
  CANR2X1 U10304 ( .A(n16842), .B(Poly10[3]), .C(Poly15[54]), .D(n16849), .Z(
        n12342) );
  CANR2X1 U10305 ( .A(n16854), .B(Poly12[32]), .C(n16839), .D(
        poly7_shifted[319]), .Z(n12341) );
  CANR2X1 U10306 ( .A(n12067), .B(poly2_shifted[17]), .C(n16864), .D(
        Poly11[67]), .Z(n12340) );
  CANR2X1 U10307 ( .A(n12071), .B(Poly5[97]), .C(n16844), .D(Poly4[39]), .Z(
        n12339) );
  CAN4X1 U10308 ( .A(n12342), .B(n12341), .C(n12340), .D(n12339), .Z(n12353)
         );
  CANR2X1 U10309 ( .A(n16840), .B(poly14_shifted[242]), .C(n16853), .D(
        Poly0[212]), .Z(n12346) );
  CANR2X1 U10310 ( .A(n12084), .B(Poly10[18]), .C(n16872), .D(
        poly0_shifted[111]), .Z(n12345) );
  CANR2X1 U10311 ( .A(n16838), .B(poly12_shifted[24]), .C(n16841), .D(
        Poly3[53]), .Z(n12344) );
  CANR2X1 U10312 ( .A(n16875), .B(poly0_shifted[146]), .C(n16862), .D(
        Poly11[49]), .Z(n12343) );
  CAN4X1 U10313 ( .A(n12346), .B(n12345), .C(n12344), .D(n12343), .Z(n12352)
         );
  CANR2X1 U10314 ( .A(n16873), .B(poly10_shifted[39]), .C(n16863), .D(
        poly14_shifted[91]), .Z(n12350) );
  CANR2X1 U10315 ( .A(n16867), .B(Poly2[54]), .C(n12872), .D(
        poly1_shifted[145]), .Z(n12349) );
  CANR2X1 U10316 ( .A(n16855), .B(Poly15[31]), .C(n16877), .D(Poly11[21]), .Z(
        n12348) );
  CANR2X1 U10317 ( .A(n16865), .B(Poly15[45]), .C(n16861), .D(Poly4[47]), .Z(
        n12347) );
  CAN4X1 U10318 ( .A(n12350), .B(n12349), .C(n12348), .D(n12347), .Z(n12351)
         );
  CND4X1 U10319 ( .A(n12354), .B(n12353), .C(n12352), .D(n12351), .Z(n12355)
         );
  CAOR2X1 U10320 ( .A(polydata[1]), .B(n17495), .C(n12355), .D(n16886), .Z(
        n8685) );
  COR3X2 U10321 ( .A(n12356), .B(n12404), .C(n18184), .Z(n14944) );
  CIVX2 U10322 ( .A(n15775), .Z(n17090) );
  CEOX1 U10323 ( .A(dataselector[62]), .B(dataselector[63]), .Z(n16407) );
  CENX1 U10324 ( .A(dataselector[59]), .B(n16407), .Z(n12357) );
  CENX1 U10325 ( .A(dataselector[6]), .B(n12357), .Z(n12358) );
  CND2X1 U10326 ( .A(n12358), .B(n17453), .Z(n12360) );
  CND2X1 U10327 ( .A(n16410), .B(dataselector[13]), .Z(n12359) );
  COND3XL U10328 ( .A(n14944), .B(n17090), .C(n12360), .D(n12359), .Z(n8782)
         );
  CND2X1 U10329 ( .A(n12017), .B(n13120), .Z(n12361) );
  CANR2X1 U10330 ( .A(n17977), .B(poly13_shifted[153]), .C(n17545), .D(
        poly13_shifted[139]), .Z(n12362) );
  COND1XL U10331 ( .A(n16605), .B(n17977), .C(n12362), .Z(n10921) );
  CEOX2 U10332 ( .A(dataselector[61]), .B(dataselector[60]), .Z(n14017) );
  CENX1 U10333 ( .A(n14017), .B(dataselector[62]), .Z(n15981) );
  CENX1 U10334 ( .A(dataselector[57]), .B(n15981), .Z(n14317) );
  CEOX1 U10335 ( .A(dataselector[59]), .B(n14317), .Z(n12363) );
  CENX1 U10336 ( .A(dataselector[56]), .B(n12363), .Z(n12366) );
  CIVX2 U10337 ( .A(n12364), .Z(n16139) );
  CANR2X1 U10338 ( .A(n16350), .B(dataselector[63]), .C(n12003), .D(n18248), 
        .Z(n12365) );
  COND1XL U10339 ( .A(n17826), .B(n12366), .C(n12365), .Z(n8732) );
  CENX1 U10340 ( .A(dataselector[59]), .B(dataselector[60]), .Z(n16409) );
  CENX1 U10341 ( .A(n18239), .B(n16409), .Z(n17828) );
  CEOXL U10342 ( .A(dataselector[62]), .B(n17828), .Z(n12367) );
  CENX1 U10343 ( .A(dataselector[44]), .B(n12367), .Z(n12370) );
  CND2XL U10344 ( .A(dataselector[51]), .B(n16350), .Z(n12369) );
  CND2XL U10345 ( .A(n18176), .B(n18248), .Z(n12368) );
  COND3XL U10346 ( .A(n12370), .B(n17744), .C(n12369), .D(n12368), .Z(n8744)
         );
  CND2X1 U10347 ( .A(n17932), .B(poly5_shifted[42]), .Z(n12372) );
  CND2XL U10348 ( .A(n17504), .B(poly5_shifted[28]), .Z(n12371) );
  COND3XL U10349 ( .A(n17930), .B(n11978), .C(n12372), .D(n12371), .Z(n11498)
         );
  CENX1 U10350 ( .A(dataselector[58]), .B(dataselector[63]), .Z(n14943) );
  CENX1 U10351 ( .A(dataselector[60]), .B(dataselector[48]), .Z(n12373) );
  CENX1 U10352 ( .A(n14943), .B(n12373), .Z(n12376) );
  CND2XL U10353 ( .A(n11999), .B(n18248), .Z(n12375) );
  CND2XL U10354 ( .A(dataselector[55]), .B(n16350), .Z(n12374) );
  COND3XL U10355 ( .A(n12376), .B(n17744), .C(n12375), .D(n12374), .Z(n8740)
         );
  CENX1 U10356 ( .A(n14017), .B(dataselector[45]), .Z(n12377) );
  CENX1 U10357 ( .A(n14943), .B(n12377), .Z(n12380) );
  CND2XL U10358 ( .A(dataselector[52]), .B(n16350), .Z(n12379) );
  CND2XL U10359 ( .A(n18082), .B(n18248), .Z(n12378) );
  COND3XL U10360 ( .A(n12380), .B(n17829), .C(n12379), .D(n12378), .Z(n8743)
         );
  CND2X1 U10361 ( .A(n12704), .B(n13136), .Z(n12382) );
  CANR2X1 U10362 ( .A(n14310), .B(Poly6[16]), .C(n17527), .D(poly6_shifted[16]), .Z(n12383) );
  COND1XL U10363 ( .A(n17062), .B(n13840), .C(n12383), .Z(n9677) );
  CEOX1 U10364 ( .A(dataselector[61]), .B(dataselector[62]), .Z(n16385) );
  CIVX1 U10365 ( .A(n16385), .Z(n12384) );
  CENX1 U10366 ( .A(n12384), .B(dataselector[58]), .Z(n12386) );
  CIVX1 U10367 ( .A(n12386), .Z(n12389) );
  COND1XL U10368 ( .A(n12386), .B(n12385), .C(n17218), .Z(n12387) );
  CMXI2X1 U10369 ( .A0(dataselector[12]), .A1(n12387), .S(n15799), .Z(n12388)
         );
  COND11XL U10370 ( .A(dataselector[5]), .B(n17829), .C(n12389), .D(n12388), 
        .Z(n8783) );
  CEOX1 U10371 ( .A(Poly4[45]), .B(Poly4[47]), .Z(n17225) );
  CENX1 U10372 ( .A(n17225), .B(n15640), .Z(n17327) );
  CENX1 U10373 ( .A(Poly4[49]), .B(Poly4[55]), .Z(n12390) );
  CENX1 U10374 ( .A(n17327), .B(n12390), .Z(n15238) );
  CENX1 U10375 ( .A(Poly4[54]), .B(Poly4[58]), .Z(n15650) );
  CENX1 U10376 ( .A(n15238), .B(n15650), .Z(n14778) );
  CIVX1 U10377 ( .A(n14778), .Z(n12392) );
  CMXI2XL U10378 ( .A0(n14361), .A1(poly4_shifted[18]), .S(n18230), .Z(n12391)
         );
  COND1XL U10379 ( .A(n17259), .B(n12392), .C(n12391), .Z(n8855) );
  COND1XL U10380 ( .A(poly5_shifted[19]), .B(n18176), .C(n18175), .Z(n12393)
         );
  CIVX1 U10381 ( .A(poly5_shifted[33]), .Z(n12584) );
  CMXI2XL U10382 ( .A0(n12393), .A1(n12584), .S(n17930), .Z(n11507) );
  COND1XL U10383 ( .A(poly5_shifted[26]), .B(n18095), .C(n18094), .Z(n12394)
         );
  CIVX1 U10384 ( .A(poly5_shifted[40]), .Z(n12669) );
  CMXI2XL U10385 ( .A0(n12394), .A1(n12669), .S(n17930), .Z(n11500) );
  CAN2X1 U10386 ( .A(n12396), .B(n12395), .Z(n13579) );
  CENX1 U10387 ( .A(Poly11[73]), .B(Poly11[81]), .Z(n17680) );
  CENX1 U10388 ( .A(n17680), .B(Poly11[65]), .Z(n12397) );
  CANR2X1 U10389 ( .A(n15843), .B(Poly11[80]), .C(n16372), .D(n12397), .Z(
        n12398) );
  COND1XL U10390 ( .A(n17062), .B(n15843), .C(n12398), .Z(n11109) );
  CIVX1 U10391 ( .A(n17757), .Z(n14754) );
  CIVXL U10392 ( .A(poly7_shifted[390]), .Z(n12399) );
  CND2IX1 U10393 ( .B(n14754), .A(n12399), .Z(n12400) );
  CND2X1 U10394 ( .A(n18117), .B(n12400), .Z(n12403) );
  CND2X1 U10395 ( .A(n12401), .B(poly7_shifted[402]), .Z(n12402) );
  COND1XL U10396 ( .A(n12403), .B(n12401), .C(n12402), .Z(n9714) );
  COND1X1 U10397 ( .A(n12405), .B(n12404), .C(n17829), .Z(n15583) );
  CANR2X1 U10398 ( .A(n17376), .B(Poly15[59]), .C(n17552), .D(
        poly15_shifted[59]), .Z(n12406) );
  COND1XL U10399 ( .A(n17741), .B(n17376), .C(n12406), .Z(n9578) );
  CND2X1 U10400 ( .A(n12157), .B(n17744), .Z(n18147) );
  CANR2X1 U10401 ( .A(n17273), .B(poly7_shifted[228]), .C(n17535), .D(
        poly7_shifted[216]), .Z(n12407) );
  COND1XL U10402 ( .A(n16179), .B(n17273), .C(n12407), .Z(n9888) );
  CANR2X1 U10403 ( .A(n18191), .B(poly1_shifted[281]), .C(n16919), .D(
        poly1_shifted[270]), .Z(n12408) );
  COND1XL U10404 ( .A(n17699), .B(n18191), .C(n12408), .Z(n9087) );
  CIVXL U10405 ( .A(Poly10[18]), .Z(n12410) );
  CND2X2 U10406 ( .A(n17558), .B(n17495), .Z(n18172) );
  COND1XL U10407 ( .A(poly10_shifted[18]), .B(n18210), .C(n18172), .Z(n12409)
         );
  CMXI2XL U10408 ( .A0(n12410), .A1(n12409), .S(n13782), .Z(n11085) );
  CIVXL U10409 ( .A(Poly10[17]), .Z(n12412) );
  COND1XL U10410 ( .A(n13522), .B(poly10_shifted[17]), .C(n18193), .Z(n12411)
         );
  CMXI2XL U10411 ( .A0(n12412), .A1(n12411), .S(n13782), .Z(n11086) );
  CIVX1 U10412 ( .A(Poly10[12]), .Z(n13759) );
  CIVX2 U10413 ( .A(Poly10[20]), .Z(n13185) );
  COND1XL U10414 ( .A(n17959), .B(n13185), .C(n17751), .Z(n12413) );
  CMXI2X1 U10415 ( .A0(n12413), .A1(n13185), .S(n13572), .Z(n12414) );
  CMXI2XL U10416 ( .A0(n12414), .A1(n13731), .S(n17411), .Z(n11071) );
  CIVX2 U10417 ( .A(n15673), .Z(n17290) );
  CEOXL U10418 ( .A(Poly10[22]), .B(Poly10[38]), .Z(n12416) );
  CANR1XL U10419 ( .A(n17290), .B(n12416), .C(n12415), .Z(n12417) );
  CIVX1 U10420 ( .A(Poly10[34]), .Z(n15955) );
  CMXI2XL U10421 ( .A0(n12417), .A1(n15955), .S(n17411), .Z(n11069) );
  CANR2X1 U10422 ( .A(n17994), .B(n16843), .C(poly13_shifted[133]), .D(n16840), 
        .Z(n12421) );
  CANR2X1 U10423 ( .A(n12067), .B(poly0_shifted[199]), .C(n16862), .D(
        Poly8[76]), .Z(n12420) );
  CANR2X1 U10424 ( .A(n16875), .B(Poly11[84]), .C(n16874), .D(
        poly0_shifted[191]), .Z(n12419) );
  CANR2X1 U10425 ( .A(n16850), .B(poly15_shifted[20]), .C(n16852), .D(
        poly9_shifted[53]), .Z(n12418) );
  CAN4X1 U10426 ( .A(n12421), .B(n12420), .C(n12419), .D(n12418), .Z(n12437)
         );
  CANR2X1 U10427 ( .A(n16839), .B(poly2_shifted[55]), .C(poly8_shifted[31]), 
        .D(n16849), .Z(n12425) );
  CANR2X1 U10428 ( .A(n16844), .B(poly1_shifted[330]), .C(n16854), .D(
        poly13_shifted[520]), .Z(n12424) );
  CANR2X1 U10429 ( .A(n12071), .B(poly15_shifted[52]), .C(n16841), .D(
        poly13_shifted[282]), .Z(n12423) );
  CANR2X1 U10430 ( .A(n16867), .B(Poly0[11]), .C(poly1_shifted[82]), .D(n16837), .Z(n12422) );
  CAN4X1 U10431 ( .A(n12425), .B(n12424), .C(n12423), .D(n12422), .Z(n12436)
         );
  CANR2X1 U10432 ( .A(n16842), .B(poly8_shifted[59]), .C(n16861), .D(
        poly10_shifted[40]), .Z(n12428) );
  CANR2X1 U10433 ( .A(n16865), .B(poly13_shifted[226]), .C(n16860), .D(
        Poly6[54]), .Z(n12427) );
  CANR2X1 U10434 ( .A(n16873), .B(poly13_shifted[86]), .C(n12872), .D(
        Poly11[23]), .Z(n12426) );
  CAN4X1 U10435 ( .A(n12429), .B(n12428), .C(n12427), .D(n12426), .Z(n12435)
         );
  CANR2X1 U10436 ( .A(n16855), .B(Poly4[19]), .C(poly8_shifted[55]), .D(n12084), .Z(n12433) );
  CANR2X1 U10437 ( .A(n16853), .B(Poly15[28]), .C(n16866), .D(
        poly1_shifted[101]), .Z(n12432) );
  CANR2X1 U10438 ( .A(n16876), .B(poly13_shifted[255]), .C(n16864), .D(
        Poly2[37]), .Z(n12431) );
  CANR2X1 U10439 ( .A(n16838), .B(Poly15[15]), .C(n16877), .D(Poly10[37]), .Z(
        n12430) );
  CAN4X1 U10440 ( .A(n12433), .B(n12432), .C(n12431), .D(n12430), .Z(n12434)
         );
  CND4X1 U10441 ( .A(n12437), .B(n12436), .C(n12435), .D(n12434), .Z(n12438)
         );
  CAOR2X1 U10442 ( .A(polydata[10]), .B(n17826), .C(n12438), .D(n16886), .Z(
        n8694) );
  CIVX3 U10443 ( .A(n17812), .Z(n15338) );
  CIVX2 U10444 ( .A(entrophy[12]), .Z(n15106) );
  CANR2X1 U10445 ( .A(n15330), .B(datain[0]), .C(entrophy[6]), .D(n11971), .Z(
        n12440) );
  CANR2XL U10446 ( .A(n17787), .B(datain[3]), .C(scrambler[28]), .D(n17495), 
        .Z(n12439) );
  COND3X1 U10447 ( .A(n15338), .B(n15106), .C(n12440), .D(n12439), .Z(n12443)
         );
  CND2X1 U10448 ( .A(n14695), .B(datain[7]), .Z(n14890) );
  CND2X1 U10449 ( .A(n15256), .B(entrophy[18]), .Z(n13949) );
  CIVX2 U10450 ( .A(entrophy[11]), .Z(n14999) );
  CNR2X1 U10451 ( .A(n14633), .B(n14999), .Z(n15159) );
  CND2X1 U10452 ( .A(n15159), .B(dataselector[25]), .Z(n14590) );
  CNR2X1 U10453 ( .A(n14981), .B(n13947), .Z(n15091) );
  CIVX2 U10454 ( .A(entrophy[24]), .Z(n14926) );
  CNR2X1 U10455 ( .A(n14473), .B(n14926), .Z(n14630) );
  CIVX2 U10456 ( .A(n15145), .Z(n15112) );
  COAN1X1 U10457 ( .A(n12441), .B(n14630), .C(n15145), .Z(n12442) );
  CNR2X1 U10458 ( .A(n12443), .B(n12442), .Z(n12466) );
  CND2X1 U10459 ( .A(n14131), .B(datain[6]), .Z(n15248) );
  COND3XL U10460 ( .A(entrophy[7]), .B(n14085), .C(n12444), .D(n14139), .Z(
        n12446) );
  CND2X2 U10461 ( .A(n14695), .B(n12216), .Z(n15108) );
  CIVX2 U10462 ( .A(n15108), .Z(n17775) );
  CANR2X1 U10463 ( .A(n17775), .B(entrophy[10]), .C(entrophy[18]), .D(n17774), 
        .Z(n12445) );
  COND4CX1 U10464 ( .A(n15248), .B(n12446), .C(n17778), .D(n12445), .Z(n12455)
         );
  CND2X1 U10465 ( .A(n14540), .B(entrophy[21]), .Z(n17760) );
  CND2X1 U10466 ( .A(n12019), .B(entrophy[10]), .Z(n12512) );
  CIVX1 U10467 ( .A(n12512), .Z(n12450) );
  CAN2X1 U10468 ( .A(n15299), .B(n14395), .Z(n12447) );
  CND2X4 U10469 ( .A(n12448), .B(n12447), .Z(n14230) );
  CIVX1 U10470 ( .A(entrophy[13]), .Z(n14225) );
  CNR2X1 U10471 ( .A(n14230), .B(n14225), .Z(n12449) );
  CIVX2 U10472 ( .A(n14640), .Z(n17792) );
  CND2X2 U10473 ( .A(n17792), .B(entrophy[9]), .Z(n14647) );
  CIVX2 U10474 ( .A(n15093), .Z(n14811) );
  CNR3X2 U10475 ( .A(n12450), .B(n12449), .C(n14811), .Z(n12452) );
  CND2X1 U10476 ( .A(n14826), .B(entrophy[17]), .Z(n14560) );
  CND2X1 U10477 ( .A(n15256), .B(entrophy[8]), .Z(n14469) );
  CAN2X1 U10478 ( .A(n14560), .B(n14469), .Z(n12451) );
  CND3X1 U10479 ( .A(n17760), .B(n12452), .C(n12451), .Z(n12453) );
  CAN2X1 U10480 ( .A(n12453), .B(n15309), .Z(n12454) );
  CNR2X1 U10481 ( .A(n12455), .B(n12454), .Z(n12465) );
  CNR2X1 U10482 ( .A(n14687), .B(n12456), .Z(n14213) );
  CIVX2 U10483 ( .A(n14213), .Z(n17807) );
  CIVX2 U10484 ( .A(entrophy[1]), .Z(n14133) );
  COR3X1 U10485 ( .A(n17807), .B(n11972), .C(n14133), .Z(n14420) );
  CND2X1 U10486 ( .A(n17776), .B(entrophy[26]), .Z(n14397) );
  CIVXL U10487 ( .A(n14397), .Z(n12457) );
  CANR2XL U10488 ( .A(n12457), .B(n12553), .C(n14695), .D(n14864), .Z(n12458)
         );
  CANR1XL U10489 ( .A(n14420), .B(n12458), .C(n15334), .Z(n12463) );
  CIVDX1 U10490 ( .A(n15200), .Z0(n12459), .Z1(n13945) );
  CNR2X1 U10491 ( .A(n12459), .B(n14871), .Z(n12501) );
  CND2X1 U10492 ( .A(n15256), .B(entrophy[5]), .Z(n14912) );
  CNR2X1 U10493 ( .A(n15218), .B(n14133), .Z(n14390) );
  CND2X1 U10494 ( .A(n11974), .B(entrophy[15]), .Z(n14947) );
  CNR2X1 U10495 ( .A(n12463), .B(n12462), .Z(n12464) );
  CND3XL U10496 ( .A(n12466), .B(n12465), .C(n12464), .Z(n8728) );
  CAN2X1 U10497 ( .A(n15206), .B(entrophy[15]), .Z(n14696) );
  CIVX2 U10498 ( .A(n14696), .Z(n15138) );
  CIVX2 U10499 ( .A(entrophy[9]), .Z(n14453) );
  CNR2X1 U10500 ( .A(n14546), .B(n14453), .Z(n15199) );
  CND2X1 U10501 ( .A(n13945), .B(entrophy[18]), .Z(n14883) );
  CND2XL U10502 ( .A(n17759), .B(entrophy[12]), .Z(n12468) );
  CND2X1 U10503 ( .A(n14695), .B(datain[0]), .Z(n15137) );
  CIVXL U10504 ( .A(n15137), .Z(n12467) );
  CNR2IX1 U10505 ( .B(n12468), .A(n12467), .Z(n12469) );
  CND2X1 U10506 ( .A(n14883), .B(n12469), .Z(n12470) );
  CNR2X1 U10507 ( .A(n15199), .B(n12470), .Z(n12471) );
  CANR11X1 U10508 ( .A(n12472), .B(n15138), .C(n12471), .D(n17763), .Z(n12478)
         );
  CND2X1 U10509 ( .A(n13945), .B(entrophy[31]), .Z(n17794) );
  CNR2X1 U10510 ( .A(n14796), .B(dataselector[25]), .Z(n15035) );
  CIVX2 U10511 ( .A(entrophy[25]), .Z(n15333) );
  CNR2X1 U10512 ( .A(n15351), .B(n15333), .Z(n15195) );
  CANR1XL U10513 ( .A(n15035), .B(entrophy[14]), .C(n15195), .Z(n12473) );
  CND2X1 U10514 ( .A(n17804), .B(n14866), .Z(n15327) );
  CANR11X1 U10515 ( .A(n17794), .B(n15208), .C(n12473), .D(n15327), .Z(n12477)
         );
  CND2X1 U10516 ( .A(n18234), .B(entrophy[27]), .Z(n15247) );
  CND2X1 U10517 ( .A(n12018), .B(n15247), .Z(n14070) );
  CNR2X1 U10518 ( .A(n14797), .B(n15302), .Z(n14593) );
  CND2X1 U10519 ( .A(n14070), .B(n14593), .Z(n12493) );
  CND2X2 U10520 ( .A(n17805), .B(n14396), .Z(n14967) );
  CND2XL U10521 ( .A(n14687), .B(n14652), .Z(n12474) );
  CNR2X1 U10522 ( .A(n14967), .B(n12474), .Z(n14880) );
  CND2XL U10523 ( .A(n14880), .B(n17804), .Z(n12475) );
  CNR2X1 U10524 ( .A(n12493), .B(n12475), .Z(n12476) );
  CNR3X1 U10525 ( .A(n12478), .B(n12477), .C(n12476), .Z(n12496) );
  COND2XL U10526 ( .A(entrophy[0]), .B(n11972), .C(n17797), .D(entrophy[22]), 
        .Z(n12480) );
  CND2XL U10527 ( .A(n14976), .B(entrophy[20]), .Z(n12479) );
  CANR4CX1 U10528 ( .A(n17807), .B(n12480), .C(n12479), .D(n12535), .Z(n12492)
         );
  CIVX2 U10529 ( .A(entrophy[4]), .Z(n14850) );
  CNR2X1 U10530 ( .A(n15334), .B(n14850), .Z(n15046) );
  CAOR2X1 U10531 ( .A(n15043), .B(n15046), .C(datain[3]), .D(n15330), .Z(
        n12491) );
  CND2X1 U10532 ( .A(n14695), .B(entrophy[12]), .Z(n14924) );
  CNR2X2 U10533 ( .A(n14928), .B(n14672), .Z(n14970) );
  CNR2X1 U10534 ( .A(n12481), .B(n14886), .Z(n12482) );
  CANR1X1 U10535 ( .A(n14970), .B(entrophy[2]), .C(n12482), .Z(n12483) );
  CND3XL U10536 ( .A(n15329), .B(n14924), .C(n12483), .Z(n12485) );
  CIVX2 U10537 ( .A(entrophy[16]), .Z(n15001) );
  CNR2X1 U10538 ( .A(n15334), .B(n15001), .Z(n15169) );
  CNR2IX1 U10539 ( .B(n15169), .A(n15335), .Z(n12484) );
  CANR1X1 U10540 ( .A(n15346), .B(n12485), .C(n12484), .Z(n12489) );
  CIVX1 U10541 ( .A(entrophy[22]), .Z(n15300) );
  CNR3X1 U10542 ( .A(n15168), .B(n15334), .C(n15300), .Z(n12487) );
  CIVX2 U10543 ( .A(datain[0]), .Z(n15352) );
  CNR2X1 U10544 ( .A(n15334), .B(n15352), .Z(n15045) );
  CNR2X1 U10545 ( .A(n12487), .B(n12486), .Z(n12488) );
  CND2X1 U10546 ( .A(n12489), .B(n12488), .Z(n12490) );
  CNR3X1 U10547 ( .A(n12492), .B(n12491), .C(n12490), .Z(n12495) );
  CND2X1 U10548 ( .A(n14131), .B(entrophy[8]), .Z(n14384) );
  CND2X1 U10549 ( .A(n14695), .B(datain[3]), .Z(n14080) );
  CND2X1 U10550 ( .A(n14384), .B(n14080), .Z(n14803) );
  CND2X1 U10551 ( .A(n14826), .B(datain[4]), .Z(n14370) );
  CND2X1 U10552 ( .A(n17759), .B(entrophy[1]), .Z(n14217) );
  CND2X1 U10553 ( .A(n15256), .B(datain[6]), .Z(n14888) );
  CNR2X1 U10554 ( .A(n12493), .B(n14545), .Z(n14078) );
  COND11X1 U10555 ( .A(n14803), .B(n14706), .C(n14078), .D(n15314), .Z(n12494)
         );
  CND2X1 U10556 ( .A(n14033), .B(entrophy[4]), .Z(n15202) );
  COND11X1 U10557 ( .A(n14561), .B(n14687), .C(n14928), .D(n15202), .Z(n12498)
         );
  COND2X1 U10558 ( .A(n14807), .B(n11970), .C(n15338), .D(n14387), .Z(n12497)
         );
  CANR1X1 U10559 ( .A(n12216), .B(n12498), .C(n12497), .Z(n12507) );
  CANR2XL U10560 ( .A(n17787), .B(entrophy[4]), .C(scrambler[23]), .D(n17259), 
        .Z(n12506) );
  CANR2X1 U10561 ( .A(n17775), .B(datain[3]), .C(entrophy[28]), .D(n17774), 
        .Z(n12505) );
  CND2X1 U10562 ( .A(n14131), .B(entrophy[0]), .Z(n15287) );
  CND2X1 U10563 ( .A(n17759), .B(datain[0]), .Z(n14579) );
  CND2X1 U10564 ( .A(n15287), .B(n14579), .Z(n13969) );
  CIVX2 U10565 ( .A(entrophy[19]), .Z(n14795) );
  CNR2X1 U10566 ( .A(n15218), .B(n14795), .Z(n14232) );
  CIVXL U10567 ( .A(n14232), .Z(n12500) );
  CND2X2 U10568 ( .A(n11969), .B(n14139), .Z(n15149) );
  CND2X1 U10569 ( .A(n17298), .B(entrophy[6]), .Z(n15211) );
  CNR3X1 U10570 ( .A(n15149), .B(n14085), .C(n15211), .Z(n17791) );
  CIVX2 U10571 ( .A(datain[1]), .Z(n14686) );
  CNR2X1 U10572 ( .A(n15283), .B(n14686), .Z(n15005) );
  CNR2X1 U10573 ( .A(n17791), .B(n15005), .Z(n12499) );
  CIVX2 U10574 ( .A(entrophy[27]), .Z(n15301) );
  CNR2X1 U10575 ( .A(n11969), .B(n15301), .Z(n14566) );
  CND2X1 U10576 ( .A(n17797), .B(n14566), .Z(n15071) );
  CND3XL U10577 ( .A(n12500), .B(n12499), .C(n15071), .Z(n12503) );
  CIVX1 U10578 ( .A(datain[3]), .Z(n15175) );
  CNR2X1 U10579 ( .A(n15351), .B(n15175), .Z(n14681) );
  CNR2X1 U10580 ( .A(n12501), .B(n14681), .Z(n14081) );
  CIVXL U10581 ( .A(n14081), .Z(n12502) );
  COND11X1 U10582 ( .A(n13969), .B(n12503), .C(n12502), .D(n15346), .Z(n12504)
         );
  CAN4X1 U10583 ( .A(n12507), .B(n12506), .C(n12505), .D(n12504), .Z(n12519)
         );
  CNR2X1 U10584 ( .A(n15283), .B(n14133), .Z(n15021) );
  CIVX2 U10585 ( .A(entrophy[31]), .Z(n14465) );
  CNR2X1 U10586 ( .A(n15351), .B(n14465), .Z(n15250) );
  CIVXL U10587 ( .A(n14370), .Z(n12509) );
  CNR2X1 U10588 ( .A(n14226), .B(n14807), .Z(n15193) );
  CND2X1 U10589 ( .A(n17759), .B(entrophy[0]), .Z(n14891) );
  CIVX2 U10590 ( .A(n14891), .Z(n13962) );
  CNR2X1 U10591 ( .A(n13958), .B(n14886), .Z(n15130) );
  CNR2X1 U10592 ( .A(n12018), .B(n15001), .Z(n12508) );
  CNR8X1 U10593 ( .A(n14232), .B(n15021), .C(n15250), .D(n12509), .E(n15193), 
        .F(n13962), .G(n15130), .H(n12508), .Z(n12517) );
  CND2XL U10594 ( .A(n17776), .B(entrophy[25]), .Z(n12511) );
  CND2X1 U10595 ( .A(n14695), .B(entrophy[17]), .Z(n15297) );
  CND2X1 U10596 ( .A(n15256), .B(entrophy[30]), .Z(n14028) );
  CND4X1 U10597 ( .A(n12511), .B(n15297), .C(n14028), .D(n12510), .Z(n12514)
         );
  CND2X1 U10598 ( .A(n14883), .B(n12512), .Z(n12513) );
  COND11X1 U10599 ( .A(n12515), .B(n12514), .C(n12513), .D(n15220), .Z(n12516)
         );
  COAN1X1 U10600 ( .A(n15112), .B(n12517), .C(n12516), .Z(n12518) );
  CND2X1 U10601 ( .A(n12519), .B(n12518), .Z(n8723) );
  CNR2X1 U10602 ( .A(n14981), .B(n14795), .Z(n14093) );
  CNR2X1 U10603 ( .A(n15218), .B(n14966), .Z(n12536) );
  CNR2X1 U10604 ( .A(n12520), .B(n15352), .Z(n15017) );
  CND2X1 U10605 ( .A(n17759), .B(entrophy[14]), .Z(n14904) );
  CND2XL U10606 ( .A(n14904), .B(n14652), .Z(n12521) );
  CNR2X1 U10607 ( .A(n15283), .B(n14465), .Z(n15205) );
  CNR2X1 U10608 ( .A(n15351), .B(n15106), .Z(n15144) );
  CND2X1 U10609 ( .A(n14695), .B(entrophy[5]), .Z(n14690) );
  CIVX2 U10610 ( .A(n15119), .Z(n14851) );
  CIVX2 U10611 ( .A(entrophy[2]), .Z(n15219) );
  CNR2X1 U10612 ( .A(n14851), .B(n15219), .Z(n15263) );
  CND2XL U10613 ( .A(n15263), .B(n17804), .Z(n12527) );
  CND2X1 U10614 ( .A(n15319), .B(datain[1]), .Z(n15063) );
  CAOR1X1 U10615 ( .A(n15063), .B(n15137), .C(n15334), .Z(n12526) );
  CND2X1 U10616 ( .A(n17804), .B(datain[5]), .Z(n14934) );
  CNR2X1 U10617 ( .A(n14473), .B(n14934), .Z(n12524) );
  CND2X1 U10618 ( .A(n15206), .B(entrophy[8]), .Z(n15344) );
  CNR2X1 U10619 ( .A(n15334), .B(n14795), .Z(n15157) );
  CANR1XL U10620 ( .A(n15157), .B(n17759), .C(n15314), .Z(n12522) );
  COND4CX1 U10621 ( .A(n15344), .B(n13946), .C(n15334), .D(n12522), .Z(n12523)
         );
  CNR2X1 U10622 ( .A(n12524), .B(n12523), .Z(n12525) );
  CND3XL U10623 ( .A(n12527), .B(n12526), .C(n12525), .Z(n12528) );
  CIVX2 U10624 ( .A(entrophy[10]), .Z(n14808) );
  CNR2X1 U10625 ( .A(n14472), .B(n14808), .Z(n14950) );
  CND2X1 U10626 ( .A(n14826), .B(datain[1]), .Z(n15268) );
  CIVX1 U10627 ( .A(n15268), .Z(n12533) );
  CIVX2 U10628 ( .A(entrophy[7]), .Z(n14567) );
  CNR2XL U10629 ( .A(n17805), .B(n14567), .Z(n12530) );
  CND2X1 U10630 ( .A(n14887), .B(n12530), .Z(n12531) );
  CND2X1 U10631 ( .A(n15256), .B(entrophy[15]), .Z(n14578) );
  CND2X1 U10632 ( .A(n15206), .B(entrophy[23]), .Z(n14824) );
  CND4X1 U10633 ( .A(n14924), .B(n12531), .C(n14578), .D(n14824), .Z(n12532)
         );
  COR3X1 U10634 ( .A(n14950), .B(n12533), .C(n12532), .Z(n12542) );
  CANR2X1 U10635 ( .A(n15249), .B(entrophy[4]), .C(n14695), .D(entrophy[20]), 
        .Z(n12538) );
  CNR2X1 U10636 ( .A(n12535), .B(dataselector[14]), .Z(n14877) );
  CANR2X1 U10637 ( .A(n12536), .B(n14877), .C(entrophy[31]), .D(n15330), .Z(
        n12537) );
  COND1X1 U10638 ( .A(n15293), .B(n12538), .C(n12537), .Z(n12541) );
  CANR3X1 U10639 ( .A(n15351), .B(n14969), .C(n17785), .D(n14686), .Z(n12539)
         );
  CAOR1XL U10640 ( .A(scrambler[8]), .B(n17826), .C(n12539), .Z(n12540) );
  CANR3X2 U10641 ( .A(n12542), .B(n15145), .C(n12541), .D(n12540), .Z(n12544)
         );
  CND2X1 U10642 ( .A(n15101), .B(dataselector[25]), .Z(n14660) );
  CIVX2 U10643 ( .A(n15354), .Z(n15332) );
  COND2X1 U10644 ( .A(n14545), .B(n14660), .C(n15332), .D(n14795), .Z(n14413)
         );
  CND2X1 U10645 ( .A(n14413), .B(n14868), .Z(n12543) );
  CND2X1 U10646 ( .A(n12019), .B(entrophy[26]), .Z(n15094) );
  COR2X1 U10647 ( .A(n15001), .B(n14472), .Z(n15143) );
  CNR2X2 U10648 ( .A(n14672), .B(n17805), .Z(n14913) );
  CND3XL U10649 ( .A(n14913), .B(n15302), .C(entrophy[21]), .Z(n14025) );
  CND4X1 U10650 ( .A(n15094), .B(n15143), .C(n13949), .D(n14025), .Z(n12548)
         );
  CIVX2 U10651 ( .A(n14967), .Z(n14670) );
  CND2X2 U10652 ( .A(n14670), .B(n18017), .Z(n14568) );
  CANR4CX1 U10653 ( .A(n14568), .B(n17785), .C(n15338), .D(n13947), .Z(n12547)
         );
  COND2X1 U10654 ( .A(n15339), .B(n15108), .C(n11970), .D(n14659), .Z(n12546)
         );
  CANR3X1 U10655 ( .A(n12216), .B(n12548), .C(n12547), .D(n12546), .Z(n12566)
         );
  CND2X1 U10656 ( .A(n14033), .B(datain[4]), .Z(n14073) );
  CIVDX1 U10657 ( .A(n15200), .Z0(n12481), .Z1(n14084) );
  CND2X1 U10658 ( .A(n14084), .B(entrophy[24]), .Z(n15190) );
  CND2X1 U10659 ( .A(n14454), .B(entrophy[13]), .Z(n15257) );
  CND2X1 U10660 ( .A(n14695), .B(entrophy[7]), .Z(n14388) );
  CND2XL U10661 ( .A(n14540), .B(entrophy[28]), .Z(n12549) );
  CND2X1 U10662 ( .A(n15256), .B(datain[3]), .Z(n17761) );
  CND2X1 U10663 ( .A(n17759), .B(entrophy[18]), .Z(n15028) );
  CND2X1 U10664 ( .A(n14680), .B(entrophy[17]), .Z(n12554) );
  CAN8X1 U10665 ( .A(n14073), .B(n15190), .C(n15257), .D(n14388), .E(n12549), 
        .F(n17761), .G(n15028), .H(n12554), .Z(n12550) );
  CNR2X1 U10666 ( .A(n12550), .B(n12055), .Z(n12558) );
  CND2XL U10667 ( .A(n15330), .B(entrophy[10]), .Z(n12551) );
  COND1XL U10668 ( .A(n14645), .B(n12552), .C(n12551), .Z(n12557) );
  CIVX2 U10669 ( .A(n14633), .Z(n15052) );
  CAN4X1 U10670 ( .A(n14693), .B(n15052), .C(dataselector[25]), .D(entrophy[1]), .Z(n12556) );
  CND2X1 U10671 ( .A(n17759), .B(entrophy[15]), .Z(n14860) );
  CND2X1 U10672 ( .A(n14695), .B(datain[4]), .Z(n15115) );
  CND2X1 U10673 ( .A(n14868), .B(n12553), .Z(n15236) );
  CANR11X1 U10674 ( .A(n14860), .B(n15115), .C(n12554), .D(n15236), .Z(n12555)
         );
  CNR4X1 U10675 ( .A(n12558), .B(n12557), .C(n12556), .D(n12555), .Z(n12565)
         );
  CND2XL U10676 ( .A(n17759), .B(entrophy[2]), .Z(n12560) );
  CIVDX1 U10677 ( .A(n12018), .Z0(n14848), .Z1(n14473) );
  CND2X2 U10678 ( .A(n14848), .B(entrophy[2]), .Z(n15227) );
  CND2X1 U10679 ( .A(n17495), .B(scrambler[12]), .Z(n12561) );
  CND2X1 U10680 ( .A(n14540), .B(datain[7]), .Z(n15150) );
  CIVDX1 U10681 ( .A(n13958), .Z0(n14131), .Z1(n14981) );
  CND2X1 U10682 ( .A(n14131), .B(entrophy[1]), .Z(n15226) );
  CND2X1 U10683 ( .A(n15256), .B(entrophy[13]), .Z(n15328) );
  CNR2X1 U10684 ( .A(n14230), .B(n14387), .Z(n14547) );
  CND2XL U10685 ( .A(n14547), .B(n14392), .Z(n12559) );
  CND2X1 U10686 ( .A(n13945), .B(datain[3]), .Z(n14925) );
  CND8X1 U10687 ( .A(n12560), .B(n15227), .C(n12561), .D(n15150), .E(n15226), 
        .F(n15328), .G(n12559), .H(n14925), .Z(n12563) );
  CND2X1 U10688 ( .A(n12563), .B(n12562), .Z(n12564) );
  CND3XL U10689 ( .A(n12566), .B(n12564), .C(n12565), .Z(n8712) );
  CND2X1 U10690 ( .A(n17538), .B(Poly6[54]), .Z(n16957) );
  CND2X1 U10691 ( .A(n12704), .B(n13145), .Z(n12914) );
  CIVX2 U10692 ( .A(n12915), .Z(n16063) );
  CIVX2 U10693 ( .A(n16959), .Z(n16961) );
  CANR2X1 U10694 ( .A(n16063), .B(Poly6[53]), .C(Poly6[43]), .D(n16961), .Z(
        n12567) );
  COAN1X1 U10695 ( .A(n12006), .B(n14166), .C(n12567), .Z(n12568) );
  COND1XL U10696 ( .A(n16957), .B(Poly6[43]), .C(n12568), .Z(n9640) );
  CND2X1 U10697 ( .A(n12704), .B(n13118), .Z(n15405) );
  CIVX1 U10698 ( .A(Poly5[112]), .Z(n12627) );
  CIVX2 U10699 ( .A(n15960), .Z(n17316) );
  CIVX2 U10700 ( .A(n15648), .Z(n17655) );
  CANR2X1 U10701 ( .A(n17655), .B(poly0_shifted[188]), .C(n15671), .D(
        poly0_shifted[206]), .Z(n12569) );
  COND1XL U10702 ( .A(n17316), .B(n11978), .C(n12569), .Z(n9389) );
  CND2X1 U10703 ( .A(n16387), .B(n17959), .Z(n18126) );
  COND1XL U10704 ( .A(poly5_shifted[34]), .B(n13428), .C(n18126), .Z(n12571)
         );
  CIVX2 U10705 ( .A(n15378), .Z(n17050) );
  CND2X1 U10706 ( .A(n17935), .B(poly5_shifted[48]), .Z(n12570) );
  COND1XL U10707 ( .A(n12571), .B(n17935), .C(n12570), .Z(n11492) );
  CND2X1 U10708 ( .A(n17607), .B(Poly5[117]), .Z(n12604) );
  COAN1XL U10709 ( .A(Poly5[95]), .B(n12604), .C(n12949), .Z(n12574) );
  CIVX1 U10710 ( .A(Poly5[117]), .Z(n15494) );
  CAN2X1 U10711 ( .A(n18234), .B(n15494), .Z(n17926) );
  CANR2X1 U10712 ( .A(n15403), .B(poly5_shifted[123]), .C(n17926), .D(
        Poly5[95]), .Z(n12573) );
  COND1XL U10713 ( .A(n12574), .B(n13904), .C(n12573), .Z(n11417) );
  CENX1 U10714 ( .A(dataselector[57]), .B(dataselector[58]), .Z(n13796) );
  CENX1 U10715 ( .A(dataselector[60]), .B(dataselector[43]), .Z(n12575) );
  CENX1 U10716 ( .A(n13796), .B(n12575), .Z(n12578) );
  CND2XL U10717 ( .A(n18210), .B(n18248), .Z(n12577) );
  CND2XL U10718 ( .A(dataselector[50]), .B(n16350), .Z(n12576) );
  COND3XL U10719 ( .A(n12578), .B(n17826), .C(n12577), .D(n12576), .Z(n8745)
         );
  CENX1 U10720 ( .A(dataselector[59]), .B(n18239), .Z(n17821) );
  CENX1 U10721 ( .A(n17821), .B(dataselector[62]), .Z(n12579) );
  CIVX1 U10722 ( .A(n12579), .Z(n12582) );
  COND1XL U10723 ( .A(n14396), .B(n12579), .C(n17753), .Z(n12580) );
  CMXI2X1 U10724 ( .A0(n12580), .A1(dataselector[54]), .S(n16350), .Z(n12581)
         );
  COND1XL U10725 ( .A(n12582), .B(n14796), .C(n12581), .Z(n8741) );
  CANR2X1 U10726 ( .A(n14310), .B(Poly6[15]), .C(n17178), .D(poly6_shifted[15]), .Z(n12583) );
  COND1XL U10727 ( .A(n17196), .B(n14310), .C(n12583), .Z(n9678) );
  COND2X1 U10728 ( .A(n17744), .B(n12584), .C(n17935), .D(n17711), .Z(n12585)
         );
  CAOR1XL U10729 ( .A(poly5_shifted[47]), .B(n15361), .C(n12585), .Z(n11493)
         );
  CEOX1 U10730 ( .A(Poly3[76]), .B(Poly3[43]), .Z(n12586) );
  CND2X1 U10731 ( .A(n17705), .B(Poly3[82]), .Z(n16728) );
  COAN1XL U10732 ( .A(n12586), .B(n16728), .C(n11997), .Z(n12588) );
  CIVDX2 U10733 ( .A(n17589), .Z0(n12616), .Z1(n17262) );
  CIVX3 U10734 ( .A(n12616), .Z(n17587) );
  CIVX1 U10735 ( .A(Poly3[82]), .Z(n18213) );
  CAN2X1 U10736 ( .A(n17317), .B(n18213), .Z(n13255) );
  CANR2X1 U10737 ( .A(n17587), .B(Poly3[57]), .C(n12586), .D(n13255), .Z(
        n12587) );
  COND1XL U10738 ( .A(n12588), .B(n17262), .C(n12587), .Z(n8883) );
  CIVXL U10739 ( .A(Poly5[91]), .Z(n12589) );
  CIVX2 U10740 ( .A(n15648), .Z(n16999) );
  CND2X1 U10741 ( .A(n16999), .B(Poly5[113]), .Z(n13410) );
  CIVX2 U10742 ( .A(n13410), .Z(n17938) );
  CIVX2 U10743 ( .A(n13354), .Z(n18189) );
  CANR1XL U10744 ( .A(n12589), .B(n17938), .C(n18189), .Z(n12591) );
  CANR2X1 U10745 ( .A(n13904), .B(poly5_shifted[119]), .C(n17940), .D(
        Poly5[91]), .Z(n12590) );
  COND1XL U10746 ( .A(n12591), .B(n12016), .C(n12590), .Z(n11421) );
  CNIVX4 U10747 ( .A(n15671), .Z(n17314) );
  CANR2X1 U10748 ( .A(n17598), .B(poly0_shifted[167]), .C(n17314), .D(
        Poly0[167]), .Z(n12592) );
  COND1XL U10749 ( .A(n17316), .B(n17718), .C(n12592), .Z(n9410) );
  CIVX2 U10750 ( .A(n14441), .Z(n17674) );
  CIVX2 U10751 ( .A(n15648), .Z(n16702) );
  CANR2X1 U10752 ( .A(n16702), .B(poly0_shifted[153]), .C(n17671), .D(
        Poly0[153]), .Z(n12593) );
  COND1XL U10753 ( .A(n17674), .B(n17123), .C(n12593), .Z(n9424) );
  CND2X1 U10754 ( .A(n12017), .B(n13126), .Z(n12594) );
  CNIVX8 U10755 ( .A(n12594), .Z(n17592) );
  CANR2X1 U10756 ( .A(n17592), .B(Poly13[280]), .C(n17655), .D(
        poly13_shifted[280]), .Z(n12595) );
  COND1XL U10757 ( .A(n16179), .B(n17592), .C(n12595), .Z(n10780) );
  CENX1 U10758 ( .A(dataselector[57]), .B(n16384), .Z(n17830) );
  CIVX1 U10759 ( .A(poly12_shifted[62]), .Z(n12603) );
  CEOXL U10760 ( .A(Poly12[126]), .B(Poly12[30]), .Z(n12601) );
  CND2IX1 U10761 ( .B(n12601), .A(n17994), .Z(n12597) );
  CND2X1 U10762 ( .A(n17699), .B(n12597), .Z(n12599) );
  CNR2IX1 U10763 ( .B(n12599), .A(n12598), .Z(n12600) );
  CANR1XL U10764 ( .A(n12601), .B(n17995), .C(n12600), .Z(n12602) );
  COND1XL U10765 ( .A(n13511), .B(n12603), .C(n12602), .Z(n10486) );
  CIVX2 U10766 ( .A(n12604), .Z(n17925) );
  CIVX1 U10767 ( .A(Poly5[82]), .Z(n12725) );
  CANR1XL U10768 ( .A(n17925), .B(n12725), .C(n12010), .Z(n12606) );
  CANR2X1 U10769 ( .A(n12016), .B(Poly5[96]), .C(Poly5[82]), .D(n17926), .Z(
        n12605) );
  COND1XL U10770 ( .A(n12606), .B(n13904), .C(n12605), .Z(n11430) );
  CIVX1 U10771 ( .A(poly5_shifted[45]), .Z(n15418) );
  CANR2X1 U10772 ( .A(n14310), .B(Poly6[3]), .C(n17634), .D(Poly6[49]), .Z(
        n12607) );
  COND1XL U10773 ( .A(n13275), .B(n13840), .C(n12607), .Z(n9690) );
  CANR2X1 U10774 ( .A(n17592), .B(poly13_shifted[281]), .C(n17655), .D(
        poly13_shifted[267]), .Z(n12608) );
  COND1XL U10775 ( .A(n16994), .B(n17592), .C(n12608), .Z(n10793) );
  CIVX2 U10776 ( .A(n15648), .Z(n17508) );
  CANR2X1 U10777 ( .A(n17508), .B(poly0_shifted[160]), .C(n17314), .D(
        Poly0[160]), .Z(n12609) );
  COND1XL U10778 ( .A(n17316), .B(n17751), .C(n12609), .Z(n9417) );
  CIVDX1 U10779 ( .A(n12968), .Z0(n14436), .Z1(n13482) );
  CND2X1 U10780 ( .A(n13482), .B(n17829), .Z(n18022) );
  COND1XL U10781 ( .A(poly13_shifted[255]), .B(n12003), .C(n18022), .Z(n12613)
         );
  CND2X1 U10782 ( .A(n12017), .B(n12610), .Z(n12611) );
  CND2X1 U10783 ( .A(n17595), .B(poly13_shifted[269]), .Z(n12612) );
  COND1XL U10784 ( .A(n12613), .B(n17595), .C(n12612), .Z(n10805) );
  CIVX2 U10785 ( .A(Poly3[79]), .Z(n18208) );
  CIVX1 U10786 ( .A(n13766), .Z(n14516) );
  CIVX2 U10787 ( .A(n12614), .Z(n13251) );
  CIVXL U10788 ( .A(poly7_shifted[102]), .Z(n12617) );
  CND2IX1 U10789 ( .B(n14754), .A(n12617), .Z(n12618) );
  CND2X1 U10790 ( .A(n18117), .B(n12618), .Z(n12620) );
  CND2X1 U10791 ( .A(n17217), .B(poly7_shifted[114]), .Z(n12619) );
  COND1XL U10792 ( .A(n12620), .B(n17217), .C(n12619), .Z(n10002) );
  CNR2X4 U10793 ( .A(n12649), .B(n18184), .Z(n14505) );
  CIVX2 U10794 ( .A(n14505), .Z(n17506) );
  CNR2X4 U10795 ( .A(n17535), .B(n14505), .Z(n17503) );
  CANR2XL U10796 ( .A(n17503), .B(poly0_shifted[20]), .C(n17215), .D(
        Poly0[204]), .Z(n12621) );
  COND1XL U10797 ( .A(n17506), .B(n16775), .C(n12621), .Z(n9575) );
  CENX1 U10798 ( .A(Poly11[74]), .B(Poly11[82]), .Z(n17675) );
  CEOX1 U10799 ( .A(Poly11[83]), .B(n17675), .Z(n15471) );
  CENX1 U10800 ( .A(Poly11[53]), .B(n15471), .Z(n12622) );
  CANR2X1 U10801 ( .A(n15843), .B(Poly11[68]), .C(n17755), .D(n12622), .Z(
        n12623) );
  COND1XL U10802 ( .A(n17423), .B(n15843), .C(n12623), .Z(n11121) );
  CANR2X1 U10803 ( .A(n17471), .B(poly7_shifted[91]), .C(n17634), .D(
        poly7_shifted[79]), .Z(n12624) );
  COND1XL U10804 ( .A(n17196), .B(n17471), .C(n12624), .Z(n10025) );
  CANR2X1 U10805 ( .A(n12625), .B(poly7_shifted[279]), .C(n17401), .D(
        poly7_shifted[267]), .Z(n12626) );
  COND1XL U10806 ( .A(n16605), .B(n12625), .C(n12626), .Z(n9837) );
  CIVXL U10807 ( .A(Poly5[118]), .Z(n15573) );
  CANR1XL U10808 ( .A(n15573), .B(n17938), .C(n18138), .Z(n12629) );
  CANR2X1 U10809 ( .A(n17930), .B(poly5_shifted[21]), .C(n17940), .D(
        Poly5[118]), .Z(n12628) );
  COND1XL U10810 ( .A(n12629), .B(n17930), .C(n12628), .Z(n11519) );
  CENX1 U10811 ( .A(Poly11[71]), .B(Poly11[79]), .Z(n17742) );
  CEOX1 U10812 ( .A(Poly11[80]), .B(n17742), .Z(n15388) );
  CENX1 U10813 ( .A(n15388), .B(Poly11[50]), .Z(n12630) );
  CANR2X1 U10814 ( .A(n15843), .B(Poly11[65]), .C(n16540), .D(n12630), .Z(
        n12631) );
  COND1XL U10815 ( .A(n17711), .B(n15843), .C(n12631), .Z(n11124) );
  CIVXL U10816 ( .A(dataselector[60]), .Z(n12634) );
  COND1XL U10817 ( .A(dataselector[60]), .B(n14652), .C(n17036), .Z(n12632) );
  CMXI2X1 U10818 ( .A0(dataselector[21]), .A1(n12632), .S(n17831), .Z(n12633)
         );
  COND1XL U10819 ( .A(n12634), .B(n14788), .C(n12633), .Z(n8774) );
  CEOX1 U10820 ( .A(Poly11[84]), .B(Poly11[76]), .Z(n17233) );
  CEOXL U10821 ( .A(Poly11[68]), .B(n17233), .Z(n12635) );
  CANR2XL U10822 ( .A(n15843), .B(Poly11[83]), .C(n17634), .D(n12635), .Z(
        n12636) );
  COND1XL U10823 ( .A(n17664), .B(n15843), .C(n12636), .Z(n11106) );
  CND2XL U10824 ( .A(n15843), .B(Poly11[84]), .Z(n12638) );
  CMXI2X1 U10825 ( .A0(n16415), .A1(n13488), .S(Poly11[69]), .Z(n12637) );
  COND3XL U10826 ( .A(n15843), .B(n16391), .C(n12638), .D(n12637), .Z(n11105)
         );
  CIVX2 U10827 ( .A(n17259), .Z(n17356) );
  COND1XL U10828 ( .A(Poly5[111]), .B(Poly5[76]), .C(n17356), .Z(n12640) );
  CMXI2XL U10829 ( .A0(n18095), .A1(Poly5[90]), .S(n17942), .Z(n12639) );
  COND4CXL U10830 ( .A(Poly5[76]), .B(Poly5[111]), .C(n12640), .D(n12639), .Z(
        n11436) );
  CIVX2 U10831 ( .A(n15673), .Z(n16695) );
  CEOXL U10832 ( .A(Poly11[80]), .B(Poly11[59]), .Z(n12641) );
  CANR2X1 U10833 ( .A(n15843), .B(Poly11[74]), .C(n16695), .D(n12641), .Z(
        n12642) );
  COND1XL U10834 ( .A(n12014), .B(n15843), .C(n12642), .Z(n11115) );
  CENX1 U10835 ( .A(Poly11[84]), .B(n17628), .Z(n13510) );
  CEOX1 U10836 ( .A(Poly11[54]), .B(n13510), .Z(n12643) );
  CANR2X1 U10837 ( .A(n15843), .B(Poly11[69]), .C(n18234), .D(n12643), .Z(
        n12644) );
  COND1XL U10838 ( .A(n11995), .B(n15843), .C(n12644), .Z(n11120) );
  CANR11XL U10839 ( .A(n17063), .B(n17628), .C(Poly11[67]), .D(n18210), .Z(
        n12647) );
  CNR2X1 U10840 ( .A(n15246), .B(Poly11[67]), .Z(n12645) );
  CANR1XL U10841 ( .A(Poly11[82]), .B(n15843), .C(n12645), .Z(n12646) );
  COND1XL U10842 ( .A(n12647), .B(n15843), .C(n12646), .Z(n11107) );
  CIVX2 U10843 ( .A(n17359), .Z(n18212) );
  COND1XL U10844 ( .A(Poly3[57]), .B(n16728), .C(n16939), .Z(n12650) );
  CANR2X1 U10845 ( .A(n12650), .B(n18212), .C(n13255), .D(Poly3[57]), .Z(
        n12651) );
  COND1XL U10846 ( .A(n12652), .B(n18212), .C(n12651), .Z(n8869) );
  CENX1 U10847 ( .A(Poly11[72]), .B(Poly11[80]), .Z(n15844) );
  CENX1 U10848 ( .A(Poly11[85]), .B(Poly11[64]), .Z(n12653) );
  CENX1 U10849 ( .A(n15844), .B(n12653), .Z(n12654) );
  CNR2XL U10850 ( .A(n12654), .B(n17959), .Z(n12655) );
  CANR1XL U10851 ( .A(Poly11[79]), .B(n15843), .C(n12655), .Z(n12656) );
  COND1XL U10852 ( .A(n17196), .B(n15843), .C(n12656), .Z(n11110) );
  CIVX2 U10853 ( .A(Poly6[55]), .Z(n13833) );
  CANR1XL U10854 ( .A(n13499), .B(n13833), .C(n18189), .Z(n12658) );
  CNR2X1 U10855 ( .A(n17495), .B(Poly6[50]), .Z(n13498) );
  CANR2X1 U10856 ( .A(n13840), .B(poly6_shifted[19]), .C(Poly6[55]), .D(n13498), .Z(n12657) );
  COND1XL U10857 ( .A(n12658), .B(n14310), .C(n12657), .Z(n9684) );
  COND1XL U10858 ( .A(Poly0[205]), .B(Poly0[8]), .C(n17705), .Z(n12660) );
  CANR2XL U10859 ( .A(n18095), .B(n14505), .C(n17503), .D(poly0_shifted[44]), 
        .Z(n12659) );
  COND4CXL U10860 ( .A(Poly0[8]), .B(Poly0[205]), .C(n12660), .D(n12659), .Z(
        n9551) );
  COND1XL U10861 ( .A(Poly0[209]), .B(Poly0[12]), .C(n18017), .Z(n12662) );
  CANR2XL U10862 ( .A(n18105), .B(n14505), .C(n17503), .D(poly0_shifted[48]), 
        .Z(n12661) );
  COND4CXL U10863 ( .A(Poly0[12]), .B(Poly0[209]), .C(n12662), .D(n12661), .Z(
        n9547) );
  CEOXL U10864 ( .A(Poly4[50]), .B(Poly4[59]), .Z(n12665) );
  CENX1 U10865 ( .A(Poly4[54]), .B(Poly4[52]), .Z(n13927) );
  CEOX2 U10866 ( .A(Poly4[58]), .B(n13927), .Z(n15186) );
  CENX2 U10867 ( .A(n15651), .B(n15186), .Z(n14614) );
  CIVX2 U10868 ( .A(n15673), .Z(n17174) );
  COND1XL U10869 ( .A(n14614), .B(n12665), .C(n17174), .Z(n12664) );
  CMXI2X1 U10870 ( .A0(n14754), .A1(poly4_shifted[23]), .S(n18230), .Z(n12663)
         );
  COND4CX1 U10871 ( .A(n12665), .B(n14614), .C(n12664), .D(n12663), .Z(n8850)
         );
  CIVX1 U10872 ( .A(n17757), .Z(n18116) );
  CND2XL U10873 ( .A(n17942), .B(Poly5[89]), .Z(n12667) );
  CND2XL U10874 ( .A(n17655), .B(poly5_shifted[89]), .Z(n12666) );
  COND3XL U10875 ( .A(n17942), .B(n11997), .C(n12667), .D(n12666), .Z(n11437)
         );
  CIVX1 U10876 ( .A(poly5_shifted[70]), .Z(n13249) );
  COND2XL U10877 ( .A(n17959), .B(n13249), .C(n17942), .D(n17757), .Z(n12668)
         );
  CAOR1XL U10878 ( .A(poly5_shifted[84]), .B(n17942), .C(n12668), .Z(n11456)
         );
  COND2XL U10879 ( .A(n17744), .B(n12669), .C(n15378), .D(n17163), .Z(n12670)
         );
  CAOR1XL U10880 ( .A(poly5_shifted[54]), .B(n17935), .C(n12670), .Z(n11486)
         );
  CIVX1 U10881 ( .A(poly5_shifted[66]), .Z(n12980) );
  COND2XL U10882 ( .A(n17959), .B(n12980), .C(n17942), .D(n16387), .Z(n12671)
         );
  CAOR1XL U10883 ( .A(poly5_shifted[80]), .B(n17942), .C(n12671), .Z(n11460)
         );
  CEOX2 U10884 ( .A(Poly4[48]), .B(Poly4[50]), .Z(n13800) );
  CENX1 U10885 ( .A(Poly4[46]), .B(n13800), .Z(n13329) );
  CENX1 U10886 ( .A(Poly4[23]), .B(n13329), .Z(n12672) );
  CENX1 U10887 ( .A(n15640), .B(n12672), .Z(n12675) );
  COND1XL U10888 ( .A(n14614), .B(n12675), .C(n16479), .Z(n12674) );
  CMXI2X1 U10889 ( .A0(n18142), .A1(Poly4[40]), .S(n12153), .Z(n12673) );
  COND4CX1 U10890 ( .A(n12675), .B(n14614), .C(n12674), .D(n12673), .Z(n8816)
         );
  CIVX1 U10891 ( .A(Poly0[206]), .Z(n12765) );
  CND2IXL U10892 ( .B(n15648), .A(n12676), .Z(n12678) );
  CANR2XL U10893 ( .A(n18099), .B(n14505), .C(n17503), .D(poly0_shifted[45]), 
        .Z(n12677) );
  COND4CXL U10894 ( .A(Poly0[9]), .B(Poly0[206]), .C(n12678), .D(n12677), .Z(
        n9550) );
  CANR2X1 U10895 ( .A(n17306), .B(Poly2[55]), .C(n17174), .D(poly2_shifted[55]), .Z(n12679) );
  COND1XL U10896 ( .A(n12000), .B(n17306), .C(n12679), .Z(n8955) );
  CIVX2 U10897 ( .A(n15648), .Z(n17266) );
  CND2X1 U10898 ( .A(poly0_shifted[114]), .B(n17266), .Z(n12682) );
  CNR2X4 U10899 ( .A(n12680), .B(n18184), .Z(n16274) );
  COND2XL U10900 ( .A(n16274), .B(Poly0[114]), .C(n15880), .D(n18210), .Z(
        n12681) );
  CND2XL U10901 ( .A(n12682), .B(n12681), .Z(n9463) );
  COND1XL U10902 ( .A(Poly7[410]), .B(Poly7[194]), .C(n16326), .Z(n12684) );
  CMXI2XL U10903 ( .A0(n18160), .A1(poly7_shifted[218]), .S(n17273), .Z(n12683) );
  COND4CXL U10904 ( .A(Poly7[194]), .B(Poly7[410]), .C(n12684), .D(n12683), 
        .Z(n9898) );
  CEOXL U10905 ( .A(Poly7[400]), .B(Poly7[184]), .Z(n12687) );
  COND1XL U10906 ( .A(Poly7[405]), .B(n12687), .C(n18017), .Z(n12686) );
  CMXI2XL U10907 ( .A0(n12004), .A1(poly7_shifted[208]), .S(n17273), .Z(n12685) );
  COND4CXL U10908 ( .A(n12687), .B(Poly7[405]), .C(n12686), .D(n12685), .Z(
        n9908) );
  CEOXL U10909 ( .A(Poly7[405]), .B(Poly7[189]), .Z(n12690) );
  COND1XL U10910 ( .A(Poly7[410]), .B(n12690), .C(n18017), .Z(n12689) );
  CMXI2XL U10911 ( .A0(n18189), .A1(poly7_shifted[213]), .S(n17273), .Z(n12688) );
  COND4CXL U10912 ( .A(n12690), .B(Poly7[410]), .C(n12689), .D(n12688), .Z(
        n9903) );
  COND1XL U10913 ( .A(Poly7[407]), .B(Poly7[191]), .C(n18017), .Z(n12692) );
  CMXI2XL U10914 ( .A0(n16381), .A1(poly7_shifted[215]), .S(n17273), .Z(n12691) );
  COND4CXL U10915 ( .A(Poly7[191]), .B(Poly7[407]), .C(n12692), .D(n12691), 
        .Z(n9901) );
  CEOXL U10916 ( .A(Poly7[409]), .B(Poly7[188]), .Z(n12695) );
  COND1XL U10917 ( .A(\dataselector_shifted[0] ), .B(n12695), .C(n17598), .Z(
        n12694) );
  CMXI2XL U10918 ( .A0(n18142), .A1(poly7_shifted[212]), .S(n17273), .Z(n12693) );
  COND4CXL U10919 ( .A(n12695), .B(\dataselector_shifted[0] ), .C(n12694), .D(
        n12693), .Z(n9904) );
  COND1XL U10920 ( .A(Poly7[409]), .B(Poly7[193]), .C(n17634), .Z(n12697) );
  CMXI2XL U10921 ( .A0(n18219), .A1(poly7_shifted[217]), .S(n17273), .Z(n12696) );
  COND4CXL U10922 ( .A(Poly7[193]), .B(Poly7[409]), .C(n12697), .D(n12696), 
        .Z(n9899) );
  COND1XL U10923 ( .A(Poly7[406]), .B(Poly7[190]), .C(n16644), .Z(n12699) );
  CMXI2XL U10924 ( .A0(n12013), .A1(poly7_shifted[214]), .S(n17273), .Z(n12698) );
  COND4CXL U10925 ( .A(Poly7[190]), .B(Poly7[406]), .C(n12699), .D(n12698), 
        .Z(n9902) );
  COND1XL U10926 ( .A(Poly7[408]), .B(Poly7[192]), .C(n17642), .Z(n12701) );
  CMXI2XL U10927 ( .A0(n13028), .A1(poly7_shifted[216]), .S(n17273), .Z(n12700) );
  COND4CXL U10928 ( .A(Poly7[192]), .B(Poly7[408]), .C(n12701), .D(n12700), 
        .Z(n9900) );
  CND2X1 U10929 ( .A(n17607), .B(Poly6[53]), .Z(n13453) );
  CIVX2 U10930 ( .A(n13452), .Z(n13689) );
  CND2XL U10931 ( .A(n13689), .B(Poly6[25]), .Z(n12702) );
  COND3XL U10932 ( .A(Poly6[25]), .B(n13453), .C(n12702), .D(n13275), .Z(
        n12703) );
  CMX2XL U10933 ( .A0(n12703), .A1(Poly6[35]), .S(n14166), .Z(n9658) );
  CND2X2 U10934 ( .A(n12704), .B(n12994), .Z(n17564) );
  CMXI2XL U10935 ( .A0(n11986), .A1(poly7_shifted[17]), .S(n17564), .Z(n12705)
         );
  CND2X1 U10936 ( .A(n17634), .B(\dataselector_shifted[0] ), .Z(n13729) );
  CND2XL U10937 ( .A(n12705), .B(n13729), .Z(n10099) );
  CIVX1 U10938 ( .A(poly0_shifted[89]), .Z(n13440) );
  COND1XL U10939 ( .A(n17959), .B(n13440), .C(n17200), .Z(n12706) );
  CMX2XL U10940 ( .A0(n12706), .A1(poly0_shifted[107]), .S(n12291), .Z(n9488)
         );
  CEOXL U10941 ( .A(Poly15[55]), .B(Poly15[56]), .Z(n12707) );
  CEOX1 U10942 ( .A(Poly15[23]), .B(n12707), .Z(n12708) );
  COAN1XL U10943 ( .A(n14525), .B(n12708), .C(n17757), .Z(n12710) );
  CIVX2 U10944 ( .A(Poly15[49]), .Z(n18050) );
  CAN2X1 U10945 ( .A(n17280), .B(n18050), .Z(n12750) );
  CANR2X1 U10946 ( .A(n17376), .B(poly15_shifted[53]), .C(n12708), .D(n12750), 
        .Z(n12709) );
  COND1XL U10947 ( .A(n12710), .B(n17376), .C(n12709), .Z(n9599) );
  CIVX2 U10948 ( .A(Poly15[58]), .Z(n12923) );
  CENX1 U10949 ( .A(Poly15[52]), .B(Poly15[26]), .Z(n12711) );
  CEOX1 U10950 ( .A(n12923), .B(n12711), .Z(n12712) );
  COAN1XL U10951 ( .A(n16555), .B(n12712), .C(n17208), .Z(n12714) );
  CIVX2 U10952 ( .A(n16558), .Z(n16562) );
  CANR2X1 U10953 ( .A(n17376), .B(poly15_shifted[56]), .C(n12712), .D(n16562), 
        .Z(n12713) );
  COND1XL U10954 ( .A(n12714), .B(n17376), .C(n12713), .Z(n9596) );
  CENX1 U10955 ( .A(Poly2[60]), .B(Poly2[67]), .Z(n17692) );
  CEOXL U10956 ( .A(n17692), .B(Poly2[20]), .Z(n12715) );
  CNR2XL U10957 ( .A(n17959), .B(n12715), .Z(n12716) );
  CANR1XL U10958 ( .A(Poly2[32]), .B(n17306), .C(n12716), .Z(n12717) );
  COND1XL U10959 ( .A(n17751), .B(n17306), .C(n12717), .Z(n8978) );
  CIVX2 U10960 ( .A(n15648), .Z(n18047) );
  CANR2X1 U10961 ( .A(n16565), .B(n18095), .C(n18047), .D(poly15_shifted[58]), 
        .Z(n12718) );
  COND1XL U10962 ( .A(n16565), .B(n12923), .C(n12718), .Z(n9579) );
  CIVXL U10963 ( .A(poly7_shifted[230]), .Z(n12719) );
  CND2IX1 U10964 ( .B(n14754), .A(n12719), .Z(n12720) );
  CND2X1 U10965 ( .A(n18117), .B(n12720), .Z(n12722) );
  CND2XL U10966 ( .A(n17574), .B(poly7_shifted[242]), .Z(n12721) );
  COND1XL U10967 ( .A(n12722), .B(n17574), .C(n12721), .Z(n9874) );
  CND2XL U10968 ( .A(n17238), .B(poly7_shifted[85]), .Z(n12724) );
  CND2XL U10969 ( .A(n17471), .B(poly7_shifted[97]), .Z(n12723) );
  COND4CXL U10970 ( .A(n12724), .B(n17036), .C(n17471), .D(n12723), .Z(n10019)
         );
  COND1XL U10971 ( .A(poly5_shifted[82]), .B(n18210), .C(n18172), .Z(n12726)
         );
  CMXI2XL U10972 ( .A0(n12726), .A1(n12725), .S(n17942), .Z(n11444) );
  COND1XL U10973 ( .A(Poly0[206]), .B(Poly0[107]), .C(n17714), .Z(n12728) );
  CANR2XL U10974 ( .A(n15880), .B(poly0_shifted[143]), .C(n18228), .D(n16274), 
        .Z(n12727) );
  COND4CXL U10975 ( .A(Poly0[107]), .B(Poly0[206]), .C(n12728), .D(n12727), 
        .Z(n9452) );
  CANR2X1 U10976 ( .A(n17376), .B(Poly15[54]), .C(n17533), .D(
        poly15_shifted[54]), .Z(n12729) );
  COND1XL U10977 ( .A(n17001), .B(n17376), .C(n12729), .Z(n9583) );
  CIVX2 U10978 ( .A(n18209), .Z(n17361) );
  CANR2X1 U10979 ( .A(n17105), .B(poly3_shifted[75]), .C(Poly3[75]), .D(n17359), .Z(n12730) );
  COND1XL U10980 ( .A(n17361), .B(n16994), .C(n12730), .Z(n8865) );
  CANR2XL U10981 ( .A(n17755), .B(poly3_shifted[78]), .C(Poly3[78]), .D(n17359), .Z(n12731) );
  COND1XL U10982 ( .A(n17361), .B(n17699), .C(n12731), .Z(n8862) );
  COND1XL U10983 ( .A(Poly0[105]), .B(Poly0[204]), .C(n17714), .Z(n12733) );
  CANR2XL U10984 ( .A(n15880), .B(poly0_shifted[141]), .C(n18099), .D(n16274), 
        .Z(n12732) );
  COND4CXL U10985 ( .A(Poly0[204]), .B(Poly0[105]), .C(n12733), .D(n12732), 
        .Z(n9454) );
  CEOXL U10986 ( .A(Poly15[54]), .B(Poly15[55]), .Z(n12734) );
  CEOX1 U10987 ( .A(Poly15[22]), .B(n12734), .Z(n12736) );
  COAN1XL U10988 ( .A(n13420), .B(n12736), .C(n11989), .Z(n12738) );
  CIVX2 U10989 ( .A(Poly15[48]), .Z(n14321) );
  CND2X1 U10990 ( .A(n16326), .B(n14321), .Z(n14323) );
  CIVX1 U10991 ( .A(n14323), .Z(n12735) );
  CANR2X1 U10992 ( .A(n17376), .B(poly15_shifted[52]), .C(n12736), .D(n12735), 
        .Z(n12737) );
  COND1XL U10993 ( .A(n12738), .B(n17376), .C(n12737), .Z(n9600) );
  CANR2X1 U10994 ( .A(n17376), .B(Poly15[52]), .C(n16427), .D(
        poly15_shifted[52]), .Z(n12739) );
  COND1XL U10995 ( .A(n17707), .B(n17376), .C(n12739), .Z(n9585) );
  CENX1 U10996 ( .A(Poly2[58]), .B(Poly2[65]), .Z(n15971) );
  CEOXL U10997 ( .A(Poly2[46]), .B(n15971), .Z(n12740) );
  CNR2XL U10998 ( .A(n17495), .B(n12740), .Z(n12741) );
  CANR1XL U10999 ( .A(Poly2[58]), .B(n17306), .C(n12741), .Z(n12742) );
  COND1XL U11000 ( .A(n17735), .B(n17306), .C(n12742), .Z(n8952) );
  CEOXL U11001 ( .A(n17692), .B(Poly2[48]), .Z(n12743) );
  CNR2XL U11002 ( .A(n17744), .B(n12743), .Z(n12744) );
  CANR1XL U11003 ( .A(Poly2[60]), .B(n17306), .C(n12744), .Z(n12745) );
  COND1XL U11004 ( .A(n11978), .B(n17306), .C(n12745), .Z(n8950) );
  CENX1 U11005 ( .A(Poly2[69]), .B(Poly2[62]), .Z(n17685) );
  CEOXL U11006 ( .A(Poly2[22]), .B(n15971), .Z(n12746) );
  CENX1 U11007 ( .A(n17685), .B(n12746), .Z(n12747) );
  CNR2XL U11008 ( .A(n12747), .B(n17959), .Z(n12748) );
  CANR1XL U11009 ( .A(Poly2[34]), .B(n17306), .C(n12748), .Z(n12749) );
  COND1XL U11010 ( .A(n16775), .B(n17306), .C(n12749), .Z(n8976) );
  CEOX1 U11011 ( .A(Poly15[17]), .B(Poly15[50]), .Z(n12751) );
  COAN1XL U11012 ( .A(n12751), .B(n14525), .C(n17751), .Z(n12753) );
  CANR2X1 U11013 ( .A(n17376), .B(Poly15[32]), .C(n12751), .D(n12750), .Z(
        n12752) );
  COND1XL U11014 ( .A(n12753), .B(n17376), .C(n12752), .Z(n9605) );
  CENX1 U11015 ( .A(Poly2[26]), .B(Poly2[66]), .Z(n12754) );
  CENX1 U11016 ( .A(n17685), .B(n12754), .Z(n12755) );
  CNR2XL U11017 ( .A(n12755), .B(n17959), .Z(n12756) );
  CANR1XL U11018 ( .A(Poly2[38]), .B(n17306), .C(n12756), .Z(n12757) );
  COND1XL U11019 ( .A(n16779), .B(n17306), .C(n12757), .Z(n8972) );
  CANR2X1 U11020 ( .A(n17306), .B(Poly2[56]), .C(n16540), .D(poly2_shifted[56]), .Z(n12758) );
  COND1XL U11021 ( .A(n17721), .B(n17306), .C(n12758), .Z(n8954) );
  CIVDX1 U11022 ( .A(n17711), .Z0(n12020), .Z1(n17697) );
  CEOXL U11023 ( .A(Poly15[50]), .B(Poly15[51]), .Z(n12759) );
  CENX1 U11024 ( .A(Poly15[18]), .B(n12759), .Z(n12760) );
  CNR2X1 U11025 ( .A(n15673), .B(n12760), .Z(n12761) );
  CANR1XL U11026 ( .A(Poly15[33]), .B(n17376), .C(n12761), .Z(n12762) );
  COND1XL U11027 ( .A(n17697), .B(n17376), .C(n12762), .Z(n9604) );
  CND2X4 U11028 ( .A(n12763), .B(n13093), .Z(n18119) );
  CND2X1 U11029 ( .A(n11981), .B(n17959), .Z(n18134) );
  CND2X1 U11030 ( .A(n12764), .B(n17829), .Z(n18159) );
  COND1XL U11031 ( .A(poly0_shifted[206]), .B(n18160), .C(n18159), .Z(n12766)
         );
  CMXI2XL U11032 ( .A0(n12766), .A1(n12765), .S(n18119), .Z(n9371) );
  COND1XL U11033 ( .A(Poly9[24]), .B(Poly9[113]), .C(n17298), .Z(n12768) );
  CMXI2XL U11034 ( .A0(n18053), .A1(poly9_shifted[46]), .S(n13351), .Z(n12767)
         );
  COND4CXL U11035 ( .A(Poly9[113]), .B(Poly9[24]), .C(n12768), .D(n12767), .Z(
        n11270) );
  COND1XL U11036 ( .A(Poly12[111]), .B(Poly12[81]), .C(n18017), .Z(n12770) );
  CMXI2XL U11037 ( .A0(poly12_shifted[113]), .A1(n14361), .S(n18001), .Z(
        n12769) );
  COND4CXL U11038 ( .A(Poly12[81]), .B(Poly12[111]), .C(n12770), .D(n12769), 
        .Z(n10435) );
  COND1XL U11039 ( .A(Poly12[122]), .B(Poly12[92]), .C(n17317), .Z(n12772) );
  CMXI2XL U11040 ( .A0(poly12_shifted[124]), .A1(n13028), .S(n18001), .Z(
        n12771) );
  COND4CXL U11041 ( .A(Poly12[92]), .B(Poly12[122]), .C(n12772), .D(n12771), 
        .Z(n10424) );
  CIVDX2 U11042 ( .A(n16994), .Z0(n16381), .Z1(n16605) );
  CND2X1 U11043 ( .A(n16605), .B(n17829), .Z(n18150) );
  CEOXL U11044 ( .A(Poly9[23]), .B(Poly9[115]), .Z(n12775) );
  COND1XL U11045 ( .A(Poly9[112]), .B(n12775), .C(n18234), .Z(n12774) );
  CMXI2XL U11046 ( .A0(n12415), .A1(poly9_shifted[45]), .S(n13351), .Z(n12773)
         );
  COND4CXL U11047 ( .A(n12775), .B(Poly9[112]), .C(n12774), .D(n12773), .Z(
        n11271) );
  CEOXL U11048 ( .A(Poly9[110]), .B(Poly9[21]), .Z(n12779) );
  COND1XL U11049 ( .A(Poly9[113]), .B(n12779), .C(n18017), .Z(n12778) );
  CIVDX2 U11050 ( .A(n12776), .Z0(n18108), .Z1(n17751) );
  CMXI2XL U11051 ( .A0(n18108), .A1(poly9_shifted[43]), .S(n13351), .Z(n12777)
         );
  COND4CXL U11052 ( .A(n12779), .B(Poly9[113]), .C(n12778), .D(n12777), .Z(
        n11273) );
  COND1XL U11053 ( .A(Poly12[126]), .B(Poly12[96]), .C(n17998), .Z(n12781) );
  CMXI2XL U11054 ( .A0(Poly12[112]), .A1(n18167), .S(n18001), .Z(n12780) );
  COND4CXL U11055 ( .A(Poly12[96]), .B(Poly12[126]), .C(n12781), .D(n12780), 
        .Z(n10420) );
  COND1XL U11056 ( .A(Poly12[95]), .B(Poly12[125]), .C(n16787), .Z(n12783) );
  CMXI2XL U11057 ( .A0(Poly12[111]), .A1(n18206), .S(n18001), .Z(n12782) );
  COND4CXL U11058 ( .A(Poly12[125]), .B(Poly12[95]), .C(n12783), .D(n12782), 
        .Z(n10421) );
  CIVXL U11059 ( .A(Poly12[121]), .Z(n12784) );
  COND1XL U11060 ( .A(Poly12[118]), .B(Poly12[88]), .C(n16702), .Z(n12786) );
  CMXI2XL U11061 ( .A0(poly12_shifted[120]), .A1(n18142), .S(n18001), .Z(
        n12785) );
  COND4CXL U11062 ( .A(Poly12[88]), .B(Poly12[118]), .C(n12786), .D(n12785), 
        .Z(n10428) );
  COND1XL U11063 ( .A(Poly12[116]), .B(Poly12[86]), .C(n18017), .Z(n12788) );
  CMXI2XL U11064 ( .A0(poly12_shifted[118]), .A1(n18116), .S(n18001), .Z(
        n12787) );
  COND4CXL U11065 ( .A(Poly12[86]), .B(Poly12[116]), .C(n12788), .D(n12787), 
        .Z(n10430) );
  COND1XL U11066 ( .A(Poly12[115]), .B(Poly12[85]), .C(n17705), .Z(n12790) );
  CMXI2XL U11067 ( .A0(poly12_shifted[117]), .A1(n11982), .S(n18001), .Z(
        n12789) );
  COND4CXL U11068 ( .A(Poly12[85]), .B(Poly12[115]), .C(n12790), .D(n12789), 
        .Z(n10431) );
  CIVX1 U11069 ( .A(Poly10[23]), .Z(n12792) );
  COND11XL U11070 ( .A(Poly10[39]), .B(n17259), .C(n12792), .D(n13275), .Z(
        n12791) );
  CANR1XL U11071 ( .A(n16091), .B(n12792), .C(n12791), .Z(n12793) );
  CIVX2 U11072 ( .A(Poly10[35]), .Z(n14354) );
  CMXI2XL U11073 ( .A0(n12793), .A1(n14354), .S(n17411), .Z(n11068) );
  CIVXL U11074 ( .A(Poly12[122]), .Z(n12795) );
  COND1XL U11075 ( .A(poly12_shifted[122]), .B(n18095), .C(n18094), .Z(n12794)
         );
  CMXI2XL U11076 ( .A0(n12795), .A1(n12794), .S(n18001), .Z(n10410) );
  CND2X1 U11077 ( .A(n17163), .B(n17495), .Z(n18141) );
  CIVXL U11078 ( .A(Poly12[126]), .Z(n12797) );
  COND1XL U11079 ( .A(poly12_shifted[126]), .B(n18105), .C(n18104), .Z(n12796)
         );
  CMXI2XL U11080 ( .A0(n12797), .A1(n12796), .S(n18001), .Z(n10406) );
  CEOXL U11081 ( .A(Poly2[54]), .B(Poly2[66]), .Z(n12798) );
  CMXI2X1 U11082 ( .A0(n17313), .A1(n13647), .S(n12798), .Z(n12800) );
  CND2X2 U11083 ( .A(n13267), .B(n12991), .Z(n17696) );
  CMXI2XL U11084 ( .A0(n12415), .A1(Poly2[66]), .S(n17696), .Z(n12799) );
  CND2XL U11085 ( .A(n12800), .B(n12799), .Z(n8944) );
  CENX1 U11086 ( .A(scrambler[30]), .B(scrambler[27]), .Z(n17891) );
  CENX1 U11087 ( .A(scrambler[25]), .B(n17891), .Z(n17911) );
  CEOX2 U11088 ( .A(scrambler[18]), .B(scrambler[17]), .Z(n17884) );
  CENX1 U11089 ( .A(scrambler[31]), .B(scrambler[29]), .Z(n17882) );
  CENX1 U11090 ( .A(scrambler[22]), .B(n17882), .Z(n17893) );
  CEOX1 U11091 ( .A(n17854), .B(n17893), .Z(n12802) );
  CEOX2 U11092 ( .A(scrambler[28]), .B(scrambler[19]), .Z(n17880) );
  CENX1 U11093 ( .A(n17880), .B(scrambler[4]), .Z(n12801) );
  CENX1 U11094 ( .A(n12802), .B(n12801), .Z(n12803) );
  CEOXL U11095 ( .A(n17911), .B(n12803), .Z(dataout[20]) );
  CIVX1 U11096 ( .A(polydata[15]), .Z(n12826) );
  CANR2X1 U11097 ( .A(n16850), .B(poly3_shifted[21]), .C(n16840), .D(
        poly7_shifted[224]), .Z(n12807) );
  CANR2X1 U11098 ( .A(n16865), .B(poly7_shifted[130]), .C(n16861), .D(
        Poly2[31]), .Z(n12806) );
  CANR2X1 U11099 ( .A(n16875), .B(poly14_shifted[75]), .C(n16855), .D(
        Poly9[94]), .Z(n12805) );
  CANR2X1 U11100 ( .A(n16842), .B(Poly9[93]), .C(n12071), .D(Poly2[21]), .Z(
        n12804) );
  CAN4X1 U11101 ( .A(n12807), .B(n12806), .C(n12805), .D(n12804), .Z(n12824)
         );
  CANR2X1 U11102 ( .A(n16849), .B(Poly0[110]), .C(n12084), .D(Poly4[51]), .Z(
        n12811) );
  CND2X1 U11103 ( .A(n17620), .B(Poly2[63]), .Z(n17368) );
  CIVX2 U11104 ( .A(n17368), .Z(n17364) );
  CANR2X1 U11105 ( .A(n17364), .B(n16838), .C(n16839), .D(poly13_shifted[220]), 
        .Z(n12810) );
  CANR2X1 U11106 ( .A(n16843), .B(poly14_shifted[73]), .C(n16864), .D(
        poly1_shifted[313]), .Z(n12809) );
  CANR2X1 U11107 ( .A(n16841), .B(poly7_shifted[234]), .C(n16872), .D(
        poly14_shifted[269]), .Z(n12808) );
  CAN4X1 U11108 ( .A(n12811), .B(n12810), .C(n12809), .D(n12808), .Z(n12823)
         );
  CANR2X1 U11109 ( .A(n12067), .B(Poly10[0]), .C(n16844), .D(poly8_shifted[78]), .Z(n12815) );
  CANR2X1 U11110 ( .A(n16873), .B(poly1_shifted[189]), .C(n16867), .D(
        Poly6[32]), .Z(n12814) );
  CANR2X1 U11111 ( .A(n16863), .B(poly11_shifted[26]), .C(n16876), .D(
        Poly12[54]), .Z(n12813) );
  CANR2X1 U11112 ( .A(n16860), .B(Poly8[3]), .C(n16854), .D(poly15_shifted[55]), .Z(n12812) );
  CAN4X1 U11113 ( .A(n12815), .B(n12814), .C(n12813), .D(n12812), .Z(n12822)
         );
  CANR2X1 U11114 ( .A(n16853), .B(poly7_shifted[79]), .C(n16862), .D(Poly9[91]), .Z(n12820) );
  CANR2X1 U11115 ( .A(n16852), .B(poly13_shifted[495]), .C(n16874), .D(
        Poly4[26]), .Z(n12819) );
  CANR2X1 U11116 ( .A(n12872), .B(Poly13[274]), .C(n16866), .D(
        poly9_shifted[91]), .Z(n12818) );
  CIVXL U11117 ( .A(n13420), .Z(n12816) );
  CANR2X1 U11118 ( .A(n16877), .B(n12816), .C(Poly2[34]), .D(n16837), .Z(
        n12817) );
  CAN4X1 U11119 ( .A(n12820), .B(n12819), .C(n12818), .D(n12817), .Z(n12821)
         );
  CAN4X1 U11120 ( .A(n12824), .B(n12823), .C(n12822), .D(n12821), .Z(n12825)
         );
  COND2X2 U11121 ( .A(n12826), .B(n16702), .C(n12825), .D(n14852), .Z(n8699)
         );
  CIVXL U11122 ( .A(polydata[4]), .Z(n12849) );
  CIVX2 U11123 ( .A(n13453), .Z(n13691) );
  CANR2X1 U11124 ( .A(n16864), .B(n13691), .C(n16840), .D(poly4_shifted[21]), 
        .Z(n12830) );
  CANR2X1 U11125 ( .A(n16860), .B(Poly11[46]), .C(n16839), .D(
        poly1_shifted[260]), .Z(n12829) );
  CANR2X1 U11126 ( .A(n16842), .B(poly7_shifted[279]), .C(poly3_shifted[77]), 
        .D(n16837), .Z(n12828) );
  CANR2X1 U11127 ( .A(n16863), .B(poly12_shifted[84]), .C(n12872), .D(
        poly3_shifted[23]), .Z(n12827) );
  CAN4X1 U11128 ( .A(n12830), .B(n12829), .C(n12828), .D(n12827), .Z(n12847)
         );
  CANR2X1 U11129 ( .A(n16844), .B(poly0_shifted[141]), .C(n16843), .D(
        poly15_shifted[15]), .Z(n12834) );
  CANR2X1 U11130 ( .A(n16855), .B(poly3_shifted[42]), .C(n16866), .D(
        Poly14[177]), .Z(n12833) );
  CANR2X1 U11131 ( .A(n16849), .B(poly7_shifted[290]), .C(n16872), .D(
        Poly10[1]), .Z(n12832) );
  CANR2X1 U11132 ( .A(n12071), .B(poly12_shifted[19]), .C(n16875), .D(
        Poly7[187]), .Z(n12831) );
  CAN4X1 U11133 ( .A(n12834), .B(n12833), .C(n12832), .D(n12831), .Z(n12846)
         );
  CANR2X1 U11134 ( .A(n16838), .B(Poly0[109]), .C(n12084), .D(
        poly1_shifted[311]), .Z(n12838) );
  CANR2X1 U11135 ( .A(n16861), .B(poly14_shifted[65]), .C(n16854), .D(
        Poly4[35]), .Z(n12837) );
  CANR2X1 U11136 ( .A(n16841), .B(Poly11[53]), .C(n16853), .D(Poly10[34]), .Z(
        n12836) );
  CANR2X1 U11137 ( .A(n16873), .B(poly15_shifted[25]), .C(n16862), .D(
        poly14_shifted[133]), .Z(n12835) );
  CAN4X1 U11138 ( .A(n12838), .B(n12837), .C(n12836), .D(n12835), .Z(n12845)
         );
  CANR2X1 U11139 ( .A(n16865), .B(poly12_shifted[90]), .C(n16874), .D(Poly6[0]), .Z(n12843) );
  CANR2X1 U11140 ( .A(n12067), .B(poly9_shifted[89]), .C(n16867), .D(
        poly12_shifted[23]), .Z(n12842) );
  CIVXL U11141 ( .A(n13371), .Z(n12839) );
  CANR2X1 U11142 ( .A(n16876), .B(n12839), .C(Poly4[33]), .D(n16852), .Z(
        n12841) );
  CANR2X1 U11143 ( .A(n16850), .B(Poly11[43]), .C(n16877), .D(
        poly3_shifted[22]), .Z(n12840) );
  CAN4X1 U11144 ( .A(n12843), .B(n12842), .C(n12841), .D(n12840), .Z(n12844)
         );
  CAN4X1 U11145 ( .A(n12847), .B(n12846), .C(n12845), .D(n12844), .Z(n12848)
         );
  COND2X2 U11146 ( .A(n12849), .B(n17613), .C(n12848), .D(n14852), .Z(n8688)
         );
  CIVXL U11147 ( .A(polydata[5]), .Z(n12871) );
  CANR2X1 U11148 ( .A(n16874), .B(poly13_shifted[493]), .C(n16866), .D(
        Poly15[21]), .Z(n12853) );
  CANR2X1 U11149 ( .A(n16838), .B(poly13_shifted[165]), .C(n16864), .D(
        poly7_shifted[349]), .Z(n12852) );
  CANR2X1 U11150 ( .A(n16855), .B(poly7_shifted[361]), .C(n16862), .D(
        Poly6[41]), .Z(n12851) );
  CANR2X1 U11151 ( .A(n16863), .B(poly15_shifted[23]), .C(n16839), .D(
        Poly11[32]), .Z(n12850) );
  CAN4X1 U11152 ( .A(n12853), .B(n12852), .C(n12851), .D(n12850), .Z(n12869)
         );
  CANR2X1 U11153 ( .A(n16865), .B(poly2_shifted[56]), .C(n16843), .D(Poly9[17]), .Z(n12857) );
  CANR2X1 U11154 ( .A(n16876), .B(poly14_shifted[169]), .C(n12872), .D(
        poly12_shifted[62]), .Z(n12856) );
  CANR2X1 U11155 ( .A(n16875), .B(Poly3[31]), .C(n12067), .D(Poly11[17]), .Z(
        n12855) );
  CANR2X1 U11156 ( .A(n16861), .B(Poly11[38]), .C(Poly2[36]), .D(n16849), .Z(
        n12854) );
  CAN4X1 U11157 ( .A(n12857), .B(n12856), .C(n12855), .D(n12854), .Z(n12868)
         );
  CANR2X1 U11158 ( .A(n16850), .B(Poly2[62]), .C(n16853), .D(
        poly1_shifted[100]), .Z(n12861) );
  CANR2X1 U11159 ( .A(n16840), .B(poly9_shifted[79]), .C(n16860), .D(Poly3[32]), .Z(n12860) );
  CANR2X1 U11160 ( .A(poly12_shifted[54]), .B(n16842), .C(Poly10[38]), .D(
        n16852), .Z(n12859) );
  CANR2X1 U11161 ( .A(n16844), .B(poly15_shifted[24]), .C(n16873), .D(
        Poly5[85]), .Z(n12858) );
  CAN4X1 U11162 ( .A(n12861), .B(n12860), .C(n12859), .D(n12858), .Z(n12867)
         );
  CANR2X1 U11163 ( .A(n16841), .B(poly5_shifted[52]), .C(poly5_shifted[24]), 
        .D(n16837), .Z(n12865) );
  CANR2X1 U11164 ( .A(n12071), .B(Poly8[74]), .C(n16854), .D(
        poly7_shifted[410]), .Z(n12864) );
  CANR2X1 U11165 ( .A(n12084), .B(Poly3[58]), .C(n16877), .D(
        poly0_shifted[194]), .Z(n12863) );
  CANR2X1 U11166 ( .A(n16867), .B(poly1_shifted[318]), .C(n16872), .D(
        Poly8[90]), .Z(n12862) );
  CAN4X1 U11167 ( .A(n12865), .B(n12864), .C(n12863), .D(n12862), .Z(n12866)
         );
  CAN4X1 U11168 ( .A(n12869), .B(n12868), .C(n12867), .D(n12866), .Z(n12870)
         );
  CIVDX1 U11169 ( .A(n14852), .Z0(n16886) );
  COND2X2 U11170 ( .A(n12871), .B(n17280), .C(n12870), .D(n14852), .Z(n8689)
         );
  CIVXL U11171 ( .A(polydata[0]), .Z(n12895) );
  CANR2X1 U11172 ( .A(n16844), .B(poly7_shifted[18]), .C(n16873), .D(
        poly3_shifted[81]), .Z(n12876) );
  CANR2X1 U11173 ( .A(n16876), .B(Poly8[1]), .C(n16860), .D(poly0_shifted[157]), .Z(n12875) );
  CANR2X1 U11174 ( .A(n12872), .B(poly5_shifted[19]), .C(n16877), .D(
        poly14_shifted[289]), .Z(n12874) );
  CANR2X1 U11175 ( .A(n16843), .B(poly1_shifted[177]), .C(poly3_shifted[27]), 
        .D(n16849), .Z(n12873) );
  CAN4X1 U11176 ( .A(n12876), .B(n12875), .C(n12874), .D(n12873), .Z(n12893)
         );
  CANR2X1 U11177 ( .A(n16840), .B(poly8_shifted[37]), .C(n16852), .D(
        poly5_shifted[25]), .Z(n12881) );
  CANR2X1 U11178 ( .A(n16838), .B(poly8_shifted[38]), .C(n16839), .D(
        poly8_shifted[35]), .Z(n12880) );
  CANR2X1 U11179 ( .A(n16842), .B(poly0_shifted[89]), .C(n16861), .D(
        poly9_shifted[52]), .Z(n12879) );
  CIVXL U11180 ( .A(n13756), .Z(n12877) );
  CANR2X1 U11181 ( .A(n12084), .B(Poly6[24]), .C(n16874), .D(n12877), .Z(
        n12878) );
  CAN4X1 U11182 ( .A(n12881), .B(n12880), .C(n12879), .D(n12878), .Z(n12892)
         );
  CANR2X1 U11183 ( .A(n16865), .B(Poly10[40]), .C(Poly0[116]), .D(n16837), .Z(
        n12885) );
  CANR2X1 U11184 ( .A(n12071), .B(Poly13[524]), .C(n12067), .D(
        poly3_shifted[20]), .Z(n12884) );
  CANR2X1 U11185 ( .A(n16863), .B(poly9_shifted[51]), .C(n16854), .D(Poly3[46]), .Z(n12883) );
  CANR2X1 U11186 ( .A(n16853), .B(poly3_shifted[17]), .C(n16862), .D(
        Poly12[90]), .Z(n12882) );
  CAN4X1 U11187 ( .A(n12885), .B(n12884), .C(n12883), .D(n12882), .Z(n12891)
         );
  CANR2X1 U11188 ( .A(n16875), .B(poly5_shifted[50]), .C(poly0_shifted[143]), 
        .D(n16850), .Z(n12889) );
  CANR2X1 U11189 ( .A(n16864), .B(Poly14[198]), .C(n16866), .D(
        poly13_shifted[233]), .Z(n12888) );
  CANR2X1 U11190 ( .A(n16841), .B(Poly15[55]), .C(n16872), .D(
        poly2_shifted[29]), .Z(n12887) );
  CANR2X1 U11191 ( .A(n16855), .B(Poly10[14]), .C(n16867), .D(
        poly8_shifted[53]), .Z(n12886) );
  CAN4X1 U11192 ( .A(n12889), .B(n12888), .C(n12887), .D(n12886), .Z(n12890)
         );
  CAN4X1 U11193 ( .A(n12893), .B(n12892), .C(n12891), .D(n12890), .Z(n12894)
         );
  COND2X2 U11194 ( .A(n12895), .B(n17094), .C(n12894), .D(n14852), .Z(n8684)
         );
  CND2X1 U11195 ( .A(n13449), .B(n17959), .Z(n18166) );
  COND1XL U11196 ( .A(poly0_shifted[208]), .B(n12381), .C(n18166), .Z(n12896)
         );
  CIVX1 U11197 ( .A(Poly0[208]), .Z(n14337) );
  CMXI2XL U11198 ( .A0(n12896), .A1(n14337), .S(n18119), .Z(n9369) );
  CND2XL U11199 ( .A(n17711), .B(n17495), .Z(n18123) );
  COND1XL U11200 ( .A(poly0_shifted[193]), .B(n12020), .C(n18123), .Z(n12898)
         );
  CND2XL U11201 ( .A(n18119), .B(poly0_shifted[211]), .Z(n12897) );
  COND1XL U11202 ( .A(n12898), .B(n18119), .C(n12897), .Z(n9384) );
  CIVX2 U11203 ( .A(n15673), .Z(n17398) );
  CANR2X1 U11204 ( .A(n15403), .B(Poly5[124]), .C(n17398), .D(
        poly5_shifted[124]), .Z(n12899) );
  COND1XL U11205 ( .A(n11978), .B(n13904), .C(n12899), .Z(n11402) );
  CANR2X1 U11206 ( .A(n12900), .B(poly13_shifted[60]), .C(n17613), .D(
        poly13_shifted[46]), .Z(n12901) );
  COND1XL U11207 ( .A(n17699), .B(n12900), .C(n12901), .Z(n11014) );
  CIVX2 U11208 ( .A(n13449), .Z(n18167) );
  COND1XL U11209 ( .A(poly0_shifted[65]), .B(n14361), .C(n18123), .Z(n12903)
         );
  CND2X1 U11210 ( .A(n12291), .B(poly0_shifted[83]), .Z(n12902) );
  COND1XL U11211 ( .A(n12903), .B(n12291), .C(n12902), .Z(n9512) );
  CANR2X1 U11212 ( .A(n18191), .B(poly1_shifted[289]), .C(n17642), .D(
        poly1_shifted[278]), .Z(n12904) );
  COND1XL U11213 ( .A(n17753), .B(n18191), .C(n12904), .Z(n9079) );
  CIVDX2 U11214 ( .A(n17050), .Z0(n17935), .Z1(n12942) );
  CIVXL U11215 ( .A(poly5_shifted[76]), .Z(n12906) );
  CIVDX1 U11216 ( .A(n17050), .Z0(n15361), .Z1(n17047) );
  CANR2XL U11217 ( .A(n17047), .B(n18105), .C(n16702), .D(poly5_shifted[62]), 
        .Z(n12905) );
  COND1XL U11218 ( .A(n12942), .B(n12906), .C(n12905), .Z(n11464) );
  CANR2X1 U11219 ( .A(n18191), .B(poly1_shifted[277]), .C(n17178), .D(
        poly1_shifted[266]), .Z(n12907) );
  COND1XL U11220 ( .A(n12014), .B(n18191), .C(n12907), .Z(n9091) );
  COND1XL U11221 ( .A(poly0_shifted[95]), .B(n12003), .C(n18022), .Z(n12909)
         );
  CND2X1 U11222 ( .A(n12291), .B(poly0_shifted[113]), .Z(n12908) );
  COND1XL U11223 ( .A(n12909), .B(n12291), .C(n12908), .Z(n9482) );
  COND1XL U11224 ( .A(poly8_shifted[31]), .B(n12003), .C(n18022), .Z(n12911)
         );
  CND2X1 U11225 ( .A(n12175), .B(poly8_shifted[45]), .Z(n12910) );
  COND1XL U11226 ( .A(n12911), .B(n12175), .C(n12910), .Z(n11370) );
  CND2X1 U11227 ( .A(n13267), .B(n13118), .Z(n12912) );
  CNIVX8 U11228 ( .A(n12912), .Z(n17610) );
  CIVX2 U11229 ( .A(n17259), .Z(n17343) );
  CANR2X1 U11230 ( .A(n17610), .B(poly1_shifted[145]), .C(n17343), .D(
        poly1_shifted[134]), .Z(n12913) );
  COND1XL U11231 ( .A(n17757), .B(n17610), .C(n12913), .Z(n9223) );
  CIVX1 U11232 ( .A(n12914), .Z(n13837) );
  CANR2XL U11233 ( .A(n12915), .B(n11999), .C(n17290), .D(poly6_shifted[55]), 
        .Z(n12916) );
  COND1XL U11234 ( .A(n13837), .B(n13833), .C(n12916), .Z(n9638) );
  CENX1 U11235 ( .A(Poly0[165]), .B(Poly0[217]), .Z(n12918) );
  COND2X1 U11236 ( .A(n15960), .B(poly0_shifted[201]), .C(n11999), .D(n17314), 
        .Z(n12917) );
  COND1XL U11237 ( .A(n12918), .B(n17744), .C(n12917), .Z(n9394) );
  CANR2X1 U11238 ( .A(n18191), .B(poly1_shifted[270]), .C(n17466), .D(
        poly1_shifted[259]), .Z(n12919) );
  COND1XL U11239 ( .A(n13275), .B(n18191), .C(n12919), .Z(n9098) );
  CIVX2 U11240 ( .A(n15648), .Z(n17238) );
  CANR2X1 U11241 ( .A(n14310), .B(Poly6[0]), .C(n17238), .D(Poly6[46]), .Z(
        n12920) );
  COND1XL U11242 ( .A(n17751), .B(n13840), .C(n12920), .Z(n9693) );
  CANR2X1 U11243 ( .A(n12192), .B(Poly1[227]), .C(n17362), .D(
        poly1_shifted[227]), .Z(n12921) );
  COND1XL U11244 ( .A(n13275), .B(n12192), .C(n12921), .Z(n9130) );
  CEOXL U11245 ( .A(Poly15[57]), .B(Poly15[51]), .Z(n12922) );
  CEOX1 U11246 ( .A(Poly15[25]), .B(n12922), .Z(n12924) );
  COAN1XL U11247 ( .A(n14515), .B(n12924), .C(n17163), .Z(n12926) );
  CAN2X1 U11248 ( .A(n17538), .B(n12923), .Z(n13037) );
  CANR2X1 U11249 ( .A(n17376), .B(poly15_shifted[55]), .C(n12924), .D(n13037), 
        .Z(n12925) );
  COND1XL U11250 ( .A(n12926), .B(n17376), .C(n12925), .Z(n9597) );
  CEOXL U11251 ( .A(Poly8[94]), .B(Poly8[15]), .Z(n12927) );
  CANR2X1 U11252 ( .A(n12175), .B(poly8_shifted[43]), .C(n18047), .D(n12927), 
        .Z(n12928) );
  COND1XL U11253 ( .A(n17185), .B(n12175), .C(n12928), .Z(n11372) );
  CANR2X1 U11254 ( .A(n12192), .B(poly1_shifted[264]), .C(n17755), .D(
        poly1_shifted[253]), .Z(n12929) );
  COND1XL U11255 ( .A(n17185), .B(n12192), .C(n12929), .Z(n9104) );
  CANR2X1 U11256 ( .A(n17610), .B(Poly1[157]), .C(n17238), .D(
        poly1_shifted[157]), .Z(n12930) );
  COND1XL U11257 ( .A(n17185), .B(n17610), .C(n12930), .Z(n9200) );
  CANR2X1 U11258 ( .A(n17094), .B(poly0_shifted[166]), .C(n15671), .D(
        Poly0[166]), .Z(n12931) );
  COND1XL U11259 ( .A(n17316), .B(n17757), .C(n12931), .Z(n9411) );
  CANR2X1 U11260 ( .A(n12932), .B(poly14_shifted[288]), .C(n17362), .D(
        poly14_shifted[272]), .Z(n12933) );
  COND1XL U11261 ( .A(n17211), .B(n12932), .C(n12933), .Z(n10133) );
  CIVXL U11262 ( .A(poly5_shifted[68]), .Z(n12935) );
  CIVX2 U11263 ( .A(n17753), .Z(n18034) );
  CANR2X1 U11264 ( .A(n17047), .B(n18034), .C(n17613), .D(poly5_shifted[54]), 
        .Z(n12934) );
  COND1XL U11265 ( .A(n12942), .B(n12935), .C(n12934), .Z(n11472) );
  CMXI2X1 U11266 ( .A0(n18053), .A1(Poly2[35]), .S(n17306), .Z(n12939) );
  CIVX2 U11267 ( .A(n12936), .Z(n17366) );
  CENX1 U11268 ( .A(Poly2[66]), .B(Poly2[59]), .Z(n17738) );
  CENX1 U11269 ( .A(Poly2[23]), .B(n17738), .Z(n12937) );
  CMXI2X1 U11270 ( .A0(n17364), .A1(n17366), .S(n12937), .Z(n12938) );
  CND2X1 U11271 ( .A(n12939), .B(n12938), .Z(n8975) );
  CIVX2 U11272 ( .A(n15673), .Z(n17099) );
  CANR2X1 U11273 ( .A(n18018), .B(poly7_shifted[22]), .C(n17099), .D(
        Poly7[409]), .Z(n12940) );
  COND1XL U11274 ( .A(n12014), .B(n18018), .C(n12940), .Z(n10094) );
  CIVX2 U11275 ( .A(n15673), .Z(n17105) );
  CANR2X1 U11276 ( .A(n18018), .B(Poly7[24]), .C(n17105), .D(poly7_shifted[24]), .Z(n12941) );
  COND1XL U11277 ( .A(n16179), .B(n18018), .C(n12941), .Z(n10080) );
  CANR2X1 U11278 ( .A(n17574), .B(Poly7[234]), .C(n17535), .D(
        poly7_shifted[234]), .Z(n12943) );
  COND1XL U11279 ( .A(n12014), .B(n17574), .C(n12943), .Z(n9870) );
  CIVX2 U11280 ( .A(n15648), .Z(n16326) );
  CANR2X1 U11281 ( .A(n18191), .B(poly1_shifted[280]), .C(n16326), .D(
        poly1_shifted[269]), .Z(n12944) );
  COND1XL U11282 ( .A(n17090), .B(n18191), .C(n12944), .Z(n9088) );
  COND1XL U11283 ( .A(poly1_shifted[127]), .B(n12003), .C(n18022), .Z(n12946)
         );
  CND2X1 U11284 ( .A(n16425), .B(poly1_shifted[138]), .Z(n12945) );
  COND1XL U11285 ( .A(n12946), .B(n16425), .C(n12945), .Z(n9230) );
  CANR2X1 U11286 ( .A(n17053), .B(Poly1[200]), .C(n17285), .D(
        poly1_shifted[200]), .Z(n12947) );
  COND1XL U11287 ( .A(n17163), .B(n17053), .C(n12947), .Z(n9157) );
  CANR2X1 U11288 ( .A(n17053), .B(Poly1[198]), .C(n17063), .D(
        poly1_shifted[198]), .Z(n12948) );
  COND1XL U11289 ( .A(n17757), .B(n17053), .C(n12948), .Z(n9159) );
  CIVDX1 U11290 ( .A(n12949), .Z0(n15775), .Z1(n17065) );
  CIVX2 U11291 ( .A(n15673), .Z(n16323) );
  CANR2X1 U11292 ( .A(n12202), .B(Poly14[205]), .C(n16323), .D(
        poly14_shifted[205]), .Z(n12950) );
  COND1XL U11293 ( .A(n17065), .B(n12202), .C(n12950), .Z(n10200) );
  CANR2X1 U11294 ( .A(n12161), .B(Poly12[88]), .C(n17072), .D(
        poly12_shifted[88]), .Z(n12951) );
  COND1XL U11295 ( .A(n16179), .B(n12161), .C(n12951), .Z(n10444) );
  CANR2X1 U11296 ( .A(n17053), .B(poly1_shifted[206]), .C(n17063), .D(
        poly1_shifted[195]), .Z(n12952) );
  COND1XL U11297 ( .A(n13275), .B(n17053), .C(n12952), .Z(n9162) );
  CIVX2 U11298 ( .A(n14159), .Z(n17502) );
  CNR2X1 U11299 ( .A(n16700), .B(n14159), .Z(n13270) );
  CNIVX4 U11300 ( .A(n13270), .Z(n17500) );
  CANR2X1 U11301 ( .A(n17500), .B(poly0_shifted[61]), .C(n17266), .D(
        poly0_shifted[43]), .Z(n12954) );
  COND1XL U11302 ( .A(n17502), .B(n16605), .C(n12954), .Z(n9534) );
  CANR2X1 U11303 ( .A(n17610), .B(poly1_shifted[147]), .C(n17965), .D(
        poly1_shifted[136]), .Z(n12955) );
  COND1XL U11304 ( .A(n17163), .B(n17610), .C(n12955), .Z(n9221) );
  CANR2XL U11305 ( .A(n12932), .B(poly14_shifted[282]), .C(n17238), .D(
        poly14_shifted[266]), .Z(n12956) );
  COND1XL U11306 ( .A(n12014), .B(n12932), .C(n12956), .Z(n10139) );
  CANR2XL U11307 ( .A(n12932), .B(poly14_shifted[285]), .C(n17285), .D(
        poly14_shifted[269]), .Z(n12957) );
  COND1XL U11308 ( .A(n17065), .B(n12932), .C(n12957), .Z(n10136) );
  CANR2XL U11309 ( .A(n12958), .B(poly14_shifted[87]), .C(n17998), .D(
        poly14_shifted[71]), .Z(n12959) );
  COND1XL U11310 ( .A(n16939), .B(n12958), .C(n12959), .Z(n10334) );
  CANR2X1 U11311 ( .A(n18198), .B(poly1_shifted[308]), .C(n18047), .D(
        poly1_shifted[297]), .Z(n12960) );
  COND1XL U11312 ( .A(n17208), .B(n18198), .C(n12960), .Z(n9060) );
  CANR2X1 U11313 ( .A(n16702), .B(poly0_shifted[191]), .C(n15671), .D(
        poly0_shifted[209]), .Z(n12961) );
  COND1XL U11314 ( .A(n17316), .B(n17188), .C(n12961), .Z(n9386) );
  CANR2X1 U11315 ( .A(n12192), .B(Poly1[234]), .C(n17099), .D(
        poly1_shifted[234]), .Z(n12962) );
  COND1XL U11316 ( .A(n12014), .B(n12192), .C(n12962), .Z(n9123) );
  CENX1 U11317 ( .A(Poly10[40]), .B(Poly10[35]), .Z(n15948) );
  CEOXL U11318 ( .A(n15948), .B(Poly10[19]), .Z(n12964) );
  CMXI2XL U11319 ( .A0(n14436), .A1(Poly10[31]), .S(n17962), .Z(n12963) );
  COND1XL U11320 ( .A(n12964), .B(n17744), .C(n12963), .Z(n11072) );
  CMXI2XL U11321 ( .A0(n12004), .A1(Poly10[4]), .S(n17962), .Z(n12965) );
  COND1XL U11322 ( .A(n17829), .B(n14354), .C(n12965), .Z(n11099) );
  CIVXL U11323 ( .A(poly10_shifted[21]), .Z(n12967) );
  CMXI2XL U11324 ( .A0(n18241), .A1(Poly10[21]), .S(n17962), .Z(n12966) );
  COND1XL U11325 ( .A(n12967), .B(n17826), .C(n12966), .Z(n11082) );
  CIVX4 U11326 ( .A(n17942), .Z(n17045) );
  CANR2X1 U11327 ( .A(n18191), .B(poly1_shifted[298]), .C(n17755), .D(
        poly1_shifted[287]), .Z(n12969) );
  COND1XL U11328 ( .A(n17188), .B(n18191), .C(n12969), .Z(n9070) );
  CIVXL U11329 ( .A(poly10_shifted[19]), .Z(n12971) );
  CMXI2XL U11330 ( .A0(n18176), .A1(Poly10[19]), .S(n17962), .Z(n12970) );
  COND1XL U11331 ( .A(n12971), .B(n17826), .C(n12970), .Z(n11084) );
  CEOXL U11332 ( .A(Poly7[402]), .B(Poly7[407]), .Z(n12972) );
  CENX1 U11333 ( .A(Poly7[186]), .B(n12972), .Z(n12973) );
  CNR2XL U11334 ( .A(n12973), .B(n17829), .Z(n12974) );
  CANR1XL U11335 ( .A(poly7_shifted[210]), .B(n17273), .C(n12974), .Z(n12975)
         );
  COND1XL U11336 ( .A(n17757), .B(n17273), .C(n12975), .Z(n9906) );
  CANR2X1 U11337 ( .A(n18018), .B(poly7_shifted[12]), .C(n17105), .D(
        Poly7[399]), .Z(n12976) );
  COND1XL U11338 ( .A(n12011), .B(n18018), .C(n12976), .Z(n10104) );
  CANR2X1 U11339 ( .A(n12977), .B(poly7_shifted[182]), .C(n17290), .D(
        poly7_shifted[170]), .Z(n12978) );
  COND1XL U11340 ( .A(n12014), .B(n12977), .C(n12978), .Z(n9934) );
  CANR2X1 U11341 ( .A(n17047), .B(n18082), .C(n16488), .D(poly5_shifted[52]), 
        .Z(n12979) );
  COND1XL U11342 ( .A(n17047), .B(n12980), .C(n12979), .Z(n11474) );
  CANR2X1 U11343 ( .A(n17376), .B(Poly15[53]), .C(n17705), .D(
        poly15_shifted[53]), .Z(n12981) );
  COND1XL U11344 ( .A(n12006), .B(n17376), .C(n12981), .Z(n9584) );
  CANR2X1 U11345 ( .A(n16425), .B(poly1_shifted[113]), .C(n17755), .D(
        poly1_shifted[102]), .Z(n12982) );
  COND1XL U11346 ( .A(n17757), .B(n16425), .C(n12982), .Z(n9255) );
  CANR2X1 U11347 ( .A(n16425), .B(poly1_shifted[115]), .C(n17538), .D(
        poly1_shifted[104]), .Z(n12983) );
  COND1XL U11348 ( .A(n17163), .B(n16425), .C(n12983), .Z(n9253) );
  CANR2X1 U11349 ( .A(n16425), .B(poly1_shifted[118]), .C(n17755), .D(
        poly1_shifted[107]), .Z(n12984) );
  COND1XL U11350 ( .A(n16605), .B(n16425), .C(n12984), .Z(n9250) );
  CANR2X1 U11351 ( .A(n17053), .B(Poly1[206]), .C(n16427), .D(
        poly1_shifted[206]), .Z(n12985) );
  COND1XL U11352 ( .A(n12764), .B(n17053), .C(n12985), .Z(n9151) );
  CANR2X1 U11353 ( .A(n12175), .B(Poly8[14]), .C(n17705), .D(poly8_shifted[14]), .Z(n12986) );
  COND1XL U11354 ( .A(n12764), .B(n12175), .C(n12986), .Z(n11387) );
  CANR2X1 U11355 ( .A(n16425), .B(poly1_shifted[121]), .C(n17620), .D(
        poly1_shifted[110]), .Z(n12987) );
  COND1XL U11356 ( .A(n17699), .B(n16425), .C(n12987), .Z(n9247) );
  CANR2X1 U11357 ( .A(n17987), .B(poly13_shifted[459]), .C(n17552), .D(
        poly13_shifted[445]), .Z(n12989) );
  COND1XL U11358 ( .A(n17185), .B(n17987), .C(n12989), .Z(n10615) );
  CANR2X1 U11359 ( .A(n17982), .B(poly13_shifted[390]), .C(n17755), .D(
        poly13_shifted[376]), .Z(n12990) );
  COND1XL U11360 ( .A(n16179), .B(n17982), .C(n12990), .Z(n10684) );
  COND1XL U11361 ( .A(poly13_shifted[495]), .B(n18206), .C(n18163), .Z(n12993)
         );
  CND2X1 U11362 ( .A(n17491), .B(poly13_shifted[509]), .Z(n12992) );
  COND1XL U11363 ( .A(n12993), .B(n17491), .C(n12992), .Z(n10565) );
  CND2X1 U11364 ( .A(n12017), .B(n12994), .Z(n12995) );
  CIVX2 U11365 ( .A(n15648), .Z(n17362) );
  CANR2X1 U11366 ( .A(n18002), .B(poly14_shifted[41]), .C(n17362), .D(
        poly14_shifted[25]), .Z(n12996) );
  COND1XL U11367 ( .A(n11997), .B(n18002), .C(n12996), .Z(n10380) );
  CANR2X1 U11368 ( .A(n12997), .B(Poly12[25]), .C(n17508), .D(
        poly12_shifted[25]), .Z(n12998) );
  COND1XL U11369 ( .A(n11997), .B(n12997), .C(n12998), .Z(n10507) );
  CANR2X1 U11370 ( .A(n18018), .B(Poly7[29]), .C(n17533), .D(poly7_shifted[29]), .Z(n12999) );
  COND1XL U11371 ( .A(n17185), .B(n18018), .C(n12999), .Z(n10075) );
  CIVX2 U11372 ( .A(n17259), .Z(n17488) );
  CANR2X1 U11373 ( .A(n18018), .B(Poly7[25]), .C(n17488), .D(poly7_shifted[25]), .Z(n13000) );
  COND1XL U11374 ( .A(n11997), .B(n18018), .C(n13000), .Z(n10079) );
  COND1XL U11375 ( .A(poly1_shifted[255]), .B(n14436), .C(n18022), .Z(n13002)
         );
  CND2X1 U11376 ( .A(n12192), .B(poly1_shifted[266]), .Z(n13001) );
  COND1XL U11377 ( .A(n13002), .B(n12192), .C(n13001), .Z(n9102) );
  CENX1 U11378 ( .A(n18245), .B(n15981), .Z(n14022) );
  CEOXL U11379 ( .A(dataselector[28]), .B(dataselector[63]), .Z(n13003) );
  CENX1 U11380 ( .A(n14022), .B(n13003), .Z(n13005) );
  CANR2X1 U11381 ( .A(n18053), .B(n18248), .C(n16350), .D(dataselector[35]), 
        .Z(n13004) );
  COND1XL U11382 ( .A(n17826), .B(n13005), .C(n13004), .Z(n8760) );
  CIVX2 U11383 ( .A(n12020), .Z(n16950) );
  CANR2X1 U11384 ( .A(n18018), .B(poly7_shifted[13]), .C(n17488), .D(
        Poly7[400]), .Z(n13006) );
  COND1XL U11385 ( .A(n16950), .B(n18018), .C(n13006), .Z(n10103) );
  CANR2X1 U11386 ( .A(n18018), .B(poly7_shifted[25]), .C(n17488), .D(
        poly7_shifted[13]), .Z(n13007) );
  COND1XL U11387 ( .A(n17065), .B(n18018), .C(n13007), .Z(n10091) );
  CANR2X1 U11388 ( .A(n18018), .B(poly7_shifted[15]), .C(n17965), .D(
        Poly7[402]), .Z(n13008) );
  COND1XL U11389 ( .A(n13275), .B(n18018), .C(n13008), .Z(n10101) );
  CANR2X1 U11390 ( .A(n17982), .B(poly13_shifted[372]), .C(n17640), .D(
        poly13_shifted[358]), .Z(n13009) );
  COND1XL U11391 ( .A(n16779), .B(n17982), .C(n13009), .Z(n10702) );
  CANR2X1 U11392 ( .A(n17987), .B(poly13_shifted[433]), .C(n17401), .D(
        poly13_shifted[419]), .Z(n13010) );
  COND1XL U11393 ( .A(n13275), .B(n17987), .C(n13010), .Z(n10641) );
  CANR2X1 U11394 ( .A(n17987), .B(poly13_shifted[452]), .C(n17755), .D(
        poly13_shifted[438]), .Z(n13011) );
  COND1XL U11395 ( .A(n17001), .B(n17987), .C(n13011), .Z(n10622) );
  CANR2X1 U11396 ( .A(n17974), .B(poly13_shifted[120]), .C(n17755), .D(
        poly13_shifted[106]), .Z(n13012) );
  COND1XL U11397 ( .A(n12014), .B(n17974), .C(n13012), .Z(n10954) );
  CANR2X1 U11398 ( .A(n17974), .B(poly13_shifted[135]), .C(n17755), .D(
        poly13_shifted[121]), .Z(n13013) );
  COND1XL U11399 ( .A(n11997), .B(n17974), .C(n13013), .Z(n10939) );
  CEOXL U11400 ( .A(Poly13[515]), .B(Poly13[156]), .Z(n13015) );
  CANR2X1 U11401 ( .A(n13014), .B(poly13_shifted[184]), .C(n17285), .D(n13015), 
        .Z(n13016) );
  COND1XL U11402 ( .A(n12014), .B(n13014), .C(n13016), .Z(n10890) );
  CANR2X1 U11403 ( .A(n13014), .B(Poly13[168]), .C(n16540), .D(
        poly13_shifted[168]), .Z(n13017) );
  COND1XL U11404 ( .A(n17163), .B(n13014), .C(n13017), .Z(n10892) );
  CANR2X1 U11405 ( .A(n13014), .B(Poly13[163]), .C(n17755), .D(
        poly13_shifted[163]), .Z(n13018) );
  COND1XL U11406 ( .A(n13275), .B(n13014), .C(n13018), .Z(n10897) );
  CANR2X1 U11407 ( .A(n17273), .B(poly7_shifted[221]), .C(n17198), .D(
        poly7_shifted[209]), .Z(n13019) );
  COND1XL U11408 ( .A(n17173), .B(n17273), .C(n13019), .Z(n9895) );
  CANR2X1 U11409 ( .A(n17273), .B(poly7_shifted[226]), .C(n17705), .D(
        poly7_shifted[214]), .Z(n13020) );
  COND1XL U11410 ( .A(n17001), .B(n17273), .C(n13020), .Z(n9890) );
  CANR4CX1 U11411 ( .A(Poly15[33]), .B(n16555), .C(n13449), .D(n17376), .Z(
        n13021) );
  CANR2X1 U11412 ( .A(n17592), .B(Poly13[270]), .C(n17545), .D(
        poly13_shifted[270]), .Z(n13023) );
  COND1XL U11413 ( .A(n17699), .B(n17592), .C(n13023), .Z(n10790) );
  CANR2X1 U11414 ( .A(n17491), .B(poly13_shifted[504]), .C(n18047), .D(
        poly13_shifted[490]), .Z(n13024) );
  COND1XL U11415 ( .A(n12014), .B(n17491), .C(n13024), .Z(n10570) );
  CANR2X1 U11416 ( .A(n17491), .B(poly13_shifted[519]), .C(n16985), .D(
        poly13_shifted[505]), .Z(n13025) );
  COND1XL U11417 ( .A(n11997), .B(n17491), .C(n13025), .Z(n10555) );
  CANR2X1 U11418 ( .A(n17491), .B(poly13_shifted[502]), .C(n16702), .D(
        poly13_shifted[488]), .Z(n13026) );
  COND1XL U11419 ( .A(n17163), .B(n17491), .C(n13026), .Z(n10572) );
  CANR2X1 U11420 ( .A(n17491), .B(poly13_shifted[497]), .C(n16372), .D(
        poly13_shifted[483]), .Z(n13027) );
  COND1XL U11421 ( .A(n13275), .B(n17491), .C(n13027), .Z(n10577) );
  CANR2X1 U11422 ( .A(n18191), .B(poly1_shifted[279]), .C(n17714), .D(
        poly1_shifted[268]), .Z(n13029) );
  COND1XL U11423 ( .A(n17087), .B(n18191), .C(n13029), .Z(n9089) );
  CIVDX2 U11424 ( .A(n13443), .Z0(n14310), .Z1(n16962) );
  CIVX1 U11425 ( .A(poly6_shifted[18]), .Z(n13032) );
  CANR4CX1 U11426 ( .A(n16957), .B(Poly6[49]), .C(n17163), .D(n13840), .Z(
        n13030) );
  CANR1XL U11427 ( .A(n16961), .B(Poly6[49]), .C(n13030), .Z(n13031) );
  COND1XL U11428 ( .A(n16962), .B(n13032), .C(n13031), .Z(n9685) );
  COND1XL U11429 ( .A(poly0_shifted[66]), .B(n12415), .C(n18126), .Z(n13034)
         );
  CND2X1 U11430 ( .A(n12291), .B(poly0_shifted[84]), .Z(n13033) );
  COND1XL U11431 ( .A(n13034), .B(n12291), .C(n13033), .Z(n9511) );
  CIVXL U11432 ( .A(Poly15[32]), .Z(n13035) );
  CANR1XL U11433 ( .A(n13036), .B(n13035), .C(n18206), .Z(n13039) );
  CANR2X1 U11434 ( .A(n17376), .B(Poly15[47]), .C(n13037), .D(Poly15[32]), .Z(
        n13038) );
  COND1XL U11435 ( .A(n13039), .B(n17376), .C(n13038), .Z(n9590) );
  CANR2X1 U11436 ( .A(n13040), .B(poly7_shifted[348]), .C(n17535), .D(
        poly7_shifted[336]), .Z(n13041) );
  COND1XL U11437 ( .A(n17211), .B(n13040), .C(n13041), .Z(n9768) );
  CANR2X1 U11438 ( .A(n18002), .B(poly14_shifted[19]), .C(n17401), .D(
        Poly14[288]), .Z(n13042) );
  COND1XL U11439 ( .A(n13275), .B(n18002), .C(n13042), .Z(n10402) );
  CAN2XL U11440 ( .A(n18017), .B(poly1_shifted[42]), .Z(n13043) );
  CANR1XL U11441 ( .A(poly1_shifted[53]), .B(n12299), .C(n13043), .Z(n13044)
         );
  COND1XL U11442 ( .A(n12014), .B(n12299), .C(n13044), .Z(n9315) );
  CANR2X1 U11443 ( .A(n12192), .B(Poly1[232]), .C(n16427), .D(
        poly1_shifted[232]), .Z(n13045) );
  COND1XL U11444 ( .A(n17163), .B(n12192), .C(n13045), .Z(n9125) );
  CANR2X1 U11445 ( .A(n12192), .B(poly1_shifted[260]), .C(n16919), .D(
        poly1_shifted[249]), .Z(n13046) );
  COND1XL U11446 ( .A(n11997), .B(n12192), .C(n13046), .Z(n9108) );
  CIVX2 U11447 ( .A(n17259), .Z(n16312) );
  CANR2X1 U11448 ( .A(n12192), .B(Poly1[235]), .C(n16312), .D(
        poly1_shifted[235]), .Z(n13047) );
  COND1XL U11449 ( .A(n16605), .B(n12192), .C(n13047), .Z(n9122) );
  CIVXL U11450 ( .A(Poly6[13]), .Z(n13050) );
  CANR4CX1 U11451 ( .A(n16957), .B(Poly6[3]), .C(n12949), .D(n13840), .Z(
        n13048) );
  CANR1XL U11452 ( .A(Poly6[3]), .B(n16961), .C(n13048), .Z(n13049) );
  COND1XL U11453 ( .A(n16962), .B(n13050), .C(n13049), .Z(n9680) );
  CND2X1 U11454 ( .A(n12949), .B(n17829), .Z(n18156) );
  CANR2X1 U11455 ( .A(n18198), .B(poly1_shifted[319]), .C(n17072), .D(
        poly1_shifted[308]), .Z(n13051) );
  COND1XL U11456 ( .A(n17707), .B(n18198), .C(n13051), .Z(n9049) );
  CANR2X1 U11457 ( .A(n17471), .B(poly7_shifted[101]), .C(n17545), .D(
        poly7_shifted[89]), .Z(n13052) );
  COND1XL U11458 ( .A(n17200), .B(n17471), .C(n13052), .Z(n10015) );
  CIVX2 U11459 ( .A(n15673), .Z(n17206) );
  CANR2X1 U11460 ( .A(n17471), .B(poly7_shifted[105]), .C(n17206), .D(
        poly7_shifted[93]), .Z(n13053) );
  COND1XL U11461 ( .A(n17185), .B(n17471), .C(n13053), .Z(n10011) );
  CIVX2 U11462 ( .A(n15673), .Z(n17203) );
  CANR2X1 U11463 ( .A(n17471), .B(poly7_shifted[86]), .C(n17203), .D(
        poly7_shifted[74]), .Z(n13054) );
  COND1XL U11464 ( .A(n12014), .B(n17471), .C(n13054), .Z(n10030) );
  CANR2X1 U11465 ( .A(n17471), .B(poly7_shifted[98]), .C(n17203), .D(
        poly7_shifted[86]), .Z(n13055) );
  COND1XL U11466 ( .A(n17001), .B(n17471), .C(n13055), .Z(n10018) );
  CIVX1 U11467 ( .A(Poly15[54]), .Z(n16742) );
  CANR4CX1 U11468 ( .A(Poly15[28]), .B(n16740), .C(n16605), .D(n17376), .Z(
        n13056) );
  CANR2X1 U11469 ( .A(n17667), .B(poly13_shifted[209]), .C(n17705), .D(
        poly13_shifted[195]), .Z(n13058) );
  COND1XL U11470 ( .A(n13275), .B(n17667), .C(n13058), .Z(n10865) );
  CANR2X1 U11471 ( .A(n17667), .B(poly13_shifted[212]), .C(n17755), .D(
        poly13_shifted[198]), .Z(n13059) );
  COND1XL U11472 ( .A(n16779), .B(n17667), .C(n13059), .Z(n10862) );
  COND1XL U11473 ( .A(n18048), .B(poly1_shifted[145]), .C(n18193), .Z(n13061)
         );
  CND2X1 U11474 ( .A(n17610), .B(poly1_shifted[156]), .Z(n13060) );
  COND1XL U11475 ( .A(n13061), .B(n17610), .C(n13060), .Z(n9212) );
  CANR2X1 U11476 ( .A(n17667), .B(poly13_shifted[214]), .C(n17072), .D(
        poly13_shifted[200]), .Z(n13062) );
  COND1XL U11477 ( .A(n17163), .B(n17667), .C(n13062), .Z(n10860) );
  CIVX2 U11478 ( .A(n15648), .Z(n17094) );
  CANR2X1 U11479 ( .A(n17667), .B(poly13_shifted[231]), .C(n17094), .D(
        poly13_shifted[217]), .Z(n13063) );
  COND1XL U11480 ( .A(n17123), .B(n17667), .C(n13063), .Z(n10843) );
  CANR2X1 U11481 ( .A(n17667), .B(poly13_shifted[230]), .C(n16702), .D(
        poly13_shifted[216]), .Z(n13064) );
  COND1XL U11482 ( .A(n16179), .B(n17667), .C(n13064), .Z(n10844) );
  CANR2X1 U11483 ( .A(n18191), .B(poly1_shifted[288]), .C(n17362), .D(
        poly1_shifted[277]), .Z(n13065) );
  COND1XL U11484 ( .A(n12006), .B(n18191), .C(n13065), .Z(n9080) );
  CANR2X1 U11485 ( .A(n12625), .B(poly7_shifted[297]), .C(n17362), .D(
        poly7_shifted[285]), .Z(n13066) );
  COND1XL U11486 ( .A(n17185), .B(n12625), .C(n13066), .Z(n9819) );
  CANR2X1 U11487 ( .A(n12625), .B(poly7_shifted[282]), .C(n16540), .D(
        poly7_shifted[270]), .Z(n13067) );
  COND1XL U11488 ( .A(n12764), .B(n12625), .C(n13067), .Z(n9834) );
  CIVX2 U11489 ( .A(n15673), .Z(n16985) );
  CANR2X1 U11490 ( .A(n12625), .B(poly7_shifted[281]), .C(n16985), .D(
        poly7_shifted[269]), .Z(n13068) );
  COND1XL U11491 ( .A(n17065), .B(n12625), .C(n13068), .Z(n9835) );
  CANR2X1 U11492 ( .A(n18191), .B(poly1_shifted[268]), .C(n16540), .D(
        poly1_shifted[257]), .Z(n13069) );
  COND1XL U11493 ( .A(n16950), .B(n18191), .C(n13069), .Z(n9100) );
  CANR2X1 U11494 ( .A(n13070), .B(poly7_shifted[143]), .C(n17535), .D(
        poly7_shifted[131]), .Z(n13071) );
  COND1XL U11495 ( .A(n13275), .B(n13070), .C(n13071), .Z(n9973) );
  CEOXL U11496 ( .A(Poly5[124]), .B(Poly5[102]), .Z(n13072) );
  CANR2X1 U11497 ( .A(n13904), .B(Poly5[116]), .C(n16326), .D(n13072), .Z(
        n13073) );
  COND1XL U11498 ( .A(n17707), .B(n13904), .C(n13073), .Z(n11410) );
  CANR2X1 U11499 ( .A(n18018), .B(Poly7[28]), .C(n16644), .D(poly7_shifted[28]), .Z(n13074) );
  COND1XL U11500 ( .A(n11978), .B(n18018), .C(n13074), .Z(n10076) );
  CIVX2 U11501 ( .A(n15673), .Z(n17288) );
  CANR2X1 U11502 ( .A(n17273), .B(poly7_shifted[232]), .C(n17288), .D(
        poly7_shifted[220]), .Z(n13075) );
  COND1XL U11503 ( .A(n11978), .B(n17273), .C(n13075), .Z(n9884) );
  CANR2X1 U11504 ( .A(n17634), .B(poly0_shifted[57]), .C(n17500), .D(
        poly0_shifted[75]), .Z(n13076) );
  COND1XL U11505 ( .A(n17502), .B(n17123), .C(n13076), .Z(n9520) );
  CANR2X1 U11506 ( .A(n12625), .B(poly7_shifted[292]), .C(n17508), .D(
        poly7_shifted[280]), .Z(n13077) );
  COND1XL U11507 ( .A(n16179), .B(n12625), .C(n13077), .Z(n9824) );
  CEOX1 U11508 ( .A(scrambler[23]), .B(scrambler[27]), .Z(n17905) );
  CEOX1 U11509 ( .A(scrambler[29]), .B(scrambler[22]), .Z(n17851) );
  CEOX1 U11510 ( .A(n17905), .B(n17851), .Z(n13079) );
  CENX1 U11511 ( .A(polydata[12]), .B(scrambler[28]), .Z(n13078) );
  CENX1 U11512 ( .A(n13079), .B(n13078), .Z(n13080) );
  CEOXL U11513 ( .A(n17884), .B(n13080), .Z(dataout[3]) );
  CANR2X1 U11514 ( .A(n17990), .B(poly13_shifted[484]), .C(n17466), .D(
        poly13_shifted[470]), .Z(n13081) );
  COND1XL U11515 ( .A(n17001), .B(n17990), .C(n13081), .Z(n10590) );
  CANR2X1 U11516 ( .A(n12299), .B(Poly1[60]), .C(n17620), .D(poly1_shifted[60]), .Z(n13082) );
  COND1XL U11517 ( .A(n11978), .B(n12299), .C(n13082), .Z(n9297) );
  CANR2X1 U11518 ( .A(n12299), .B(poly1_shifted[54]), .C(n17072), .D(
        poly1_shifted[43]), .Z(n13083) );
  COND1XL U11519 ( .A(n16605), .B(n12299), .C(n13083), .Z(n9314) );
  CANR2X1 U11520 ( .A(n17990), .B(poly13_shifted[469]), .C(n17620), .D(
        poly13_shifted[455]), .Z(n13084) );
  COND1XL U11521 ( .A(n16939), .B(n17990), .C(n13084), .Z(n10605) );
  CANR2X1 U11522 ( .A(n17595), .B(poly13_shifted[262]), .C(n17755), .D(
        poly13_shifted[248]), .Z(n13085) );
  COND1XL U11523 ( .A(n16179), .B(n17595), .C(n13085), .Z(n10812) );
  CANR2X1 U11524 ( .A(n17595), .B(poly13_shifted[267]), .C(n17266), .D(
        poly13_shifted[253]), .Z(n13086) );
  COND1XL U11525 ( .A(n17185), .B(n17595), .C(n13086), .Z(n10807) );
  CANR2X1 U11526 ( .A(n12625), .B(poly7_shifted[293]), .C(n16985), .D(
        poly7_shifted[281]), .Z(n13087) );
  COND1XL U11527 ( .A(n17123), .B(n12625), .C(n13087), .Z(n9823) );
  CANR2X1 U11528 ( .A(n17332), .B(poly1_shifted[341]), .C(n17504), .D(
        poly1_shifted[330]), .Z(n13088) );
  COND1XL U11529 ( .A(n12014), .B(n17332), .C(n13088), .Z(n9027) );
  COND1XL U11530 ( .A(poly14_shifted[65]), .B(n13812), .C(n18123), .Z(n13090)
         );
  CND2X1 U11531 ( .A(n12958), .B(poly14_shifted[81]), .Z(n13089) );
  COND1XL U11532 ( .A(n13090), .B(n12958), .C(n13089), .Z(n10340) );
  CANR2X1 U11533 ( .A(n17990), .B(poly13_shifted[470]), .C(n17535), .D(
        poly13_shifted[456]), .Z(n13091) );
  COND1XL U11534 ( .A(n17163), .B(n17990), .C(n13091), .Z(n10604) );
  CANR2X1 U11535 ( .A(n17705), .B(poly0_shifted[139]), .C(poly0_shifted[157]), 
        .D(n17671), .Z(n13092) );
  COND1XL U11536 ( .A(n17674), .B(n16605), .C(n13092), .Z(n9438) );
  CND2X4 U11537 ( .A(n12017), .B(n13093), .Z(n17043) );
  CEOXL U11538 ( .A(Poly13[394]), .B(Poly13[521]), .Z(n13094) );
  CANR2X1 U11539 ( .A(n17043), .B(poly13_shifted[422]), .C(n16702), .D(n13094), 
        .Z(n13095) );
  COND1XL U11540 ( .A(n16179), .B(n17043), .C(n13095), .Z(n10652) );
  CANR2X1 U11541 ( .A(n17043), .B(Poly13[399]), .C(poly13_shifted[399]), .D(
        n18017), .Z(n13096) );
  COND1XL U11542 ( .A(n17196), .B(n17043), .C(n13096), .Z(n10661) );
  CANR2X1 U11543 ( .A(n17043), .B(Poly13[390]), .C(n17755), .D(
        poly13_shifted[390]), .Z(n13097) );
  COND1XL U11544 ( .A(n16779), .B(n17043), .C(n13097), .Z(n10670) );
  COND1XL U11545 ( .A(poly13_shifted[133]), .B(n11992), .C(n18134), .Z(n13099)
         );
  CND2X1 U11546 ( .A(n17977), .B(poly13_shifted[147]), .Z(n13098) );
  COND1XL U11547 ( .A(n13099), .B(n17977), .C(n13098), .Z(n10927) );
  CANR2X1 U11548 ( .A(n18028), .B(poly7_shifted[315]), .C(n17538), .D(
        poly7_shifted[303]), .Z(n13101) );
  COND1XL U11549 ( .A(n17196), .B(n18028), .C(n13101), .Z(n9801) );
  CANR2X1 U11550 ( .A(n18028), .B(poly7_shifted[300]), .C(n17535), .D(
        poly7_shifted[288]), .Z(n13102) );
  COND1XL U11551 ( .A(n12011), .B(n18028), .C(n13102), .Z(n9816) );
  CANR2X1 U11552 ( .A(n18028), .B(poly7_shifted[303]), .C(n17466), .D(
        poly7_shifted[291]), .Z(n13103) );
  COND1XL U11553 ( .A(n13275), .B(n18028), .C(n13103), .Z(n9813) );
  CANR2X1 U11554 ( .A(n18028), .B(poly7_shifted[314]), .C(n17535), .D(
        poly7_shifted[302]), .Z(n13104) );
  COND1XL U11555 ( .A(n12764), .B(n18028), .C(n13104), .Z(n9802) );
  CANR2X1 U11556 ( .A(n18028), .B(poly7_shifted[309]), .C(n17642), .D(
        poly7_shifted[297]), .Z(n13105) );
  COND1XL U11557 ( .A(n17208), .B(n18028), .C(n13105), .Z(n9807) );
  CIVX2 U11558 ( .A(n17259), .Z(n17295) );
  CANR2X1 U11559 ( .A(n18028), .B(poly7_shifted[310]), .C(n17295), .D(
        poly7_shifted[298]), .Z(n13106) );
  COND1XL U11560 ( .A(n12014), .B(n18028), .C(n13106), .Z(n9806) );
  CANR2X1 U11561 ( .A(n18028), .B(poly7_shifted[329]), .C(n17136), .D(
        poly7_shifted[317]), .Z(n13107) );
  COND1XL U11562 ( .A(n17185), .B(n18028), .C(n13107), .Z(n9787) );
  CANR2X1 U11563 ( .A(n17714), .B(poly3_shifted[77]), .C(Poly3[77]), .D(n17359), .Z(n13108) );
  COND1XL U11564 ( .A(n17361), .B(n17065), .C(n13108), .Z(n8863) );
  CANR2X1 U11565 ( .A(n17705), .B(poly0_shifted[142]), .C(n17671), .D(
        poly0_shifted[160]), .Z(n13109) );
  COND1XL U11566 ( .A(n17674), .B(n17699), .C(n13109), .Z(n9435) );
  CEOXL U11567 ( .A(Poly7[187]), .B(Poly7[403]), .Z(n13110) );
  CENX1 U11568 ( .A(Poly7[408]), .B(n13110), .Z(n13111) );
  CNR2XL U11569 ( .A(n13111), .B(n17259), .Z(n13112) );
  CANR1XL U11570 ( .A(poly7_shifted[211]), .B(n17273), .C(n13112), .Z(n13113)
         );
  COND1XL U11571 ( .A(n16939), .B(n17273), .C(n13113), .Z(n9905) );
  CANR2X1 U11572 ( .A(n12202), .B(Poly14[199]), .C(n17965), .D(
        poly14_shifted[199]), .Z(n13114) );
  COND1XL U11573 ( .A(n16939), .B(n12202), .C(n13114), .Z(n10206) );
  CANR2X1 U11574 ( .A(n17332), .B(poly1_shifted[338]), .C(n17620), .D(
        poly1_shifted[327]), .Z(n13115) );
  COND1XL U11575 ( .A(n16939), .B(n17332), .C(n13115), .Z(n9030) );
  CANR2X1 U11576 ( .A(n12625), .B(poly7_shifted[275]), .C(n16312), .D(
        poly7_shifted[263]), .Z(n13116) );
  COND1XL U11577 ( .A(n16939), .B(n12625), .C(n13116), .Z(n9841) );
  CND2X2 U11578 ( .A(n13878), .B(n13136), .Z(n17444) );
  CANR2XL U11579 ( .A(n17444), .B(Poly14[295]), .C(n17998), .D(
        poly14_shifted[295]), .Z(n13117) );
  COND1XL U11580 ( .A(n16939), .B(n17444), .C(n13117), .Z(n10110) );
  CANR2X1 U11581 ( .A(n12008), .B(poly14_shifted[151]), .C(n17705), .D(
        poly14_shifted[135]), .Z(n13119) );
  COND1XL U11582 ( .A(n16939), .B(n12008), .C(n13119), .Z(n10270) );
  CANR2X1 U11583 ( .A(n12009), .B(poly14_shifted[119]), .C(n17504), .D(
        poly14_shifted[103]), .Z(n13121) );
  COND1XL U11584 ( .A(n16939), .B(n12009), .C(n13121), .Z(n10302) );
  CANR2X1 U11585 ( .A(n13070), .B(poly7_shifted[147]), .C(n17063), .D(
        poly7_shifted[135]), .Z(n13122) );
  COND1XL U11586 ( .A(n16939), .B(n13070), .C(n13122), .Z(n9969) );
  CIVX2 U11587 ( .A(n15648), .Z(n17072) );
  CANR2X1 U11588 ( .A(n13124), .B(poly13_shifted[21]), .C(n17072), .D(
        Poly13[521]), .Z(n13125) );
  COND1XL U11589 ( .A(n16939), .B(n13124), .C(n13125), .Z(n11053) );
  CANR2X1 U11590 ( .A(n16694), .B(poly14_shifted[247]), .C(n17266), .D(
        poly14_shifted[231]), .Z(n13127) );
  COND1XL U11591 ( .A(n16939), .B(n16694), .C(n13127), .Z(n10174) );
  CANR2X1 U11592 ( .A(n13129), .B(Poly14[167]), .C(n17198), .D(
        poly14_shifted[167]), .Z(n13130) );
  COND1XL U11593 ( .A(n16939), .B(n13129), .C(n13130), .Z(n10238) );
  CANR2X1 U11594 ( .A(n17977), .B(poly13_shifted[149]), .C(n17755), .D(
        poly13_shifted[135]), .Z(n13131) );
  COND1XL U11595 ( .A(n16939), .B(n17977), .C(n13131), .Z(n10925) );
  CANR2X1 U11596 ( .A(n12977), .B(poly7_shifted[179]), .C(n17245), .D(
        poly7_shifted[167]), .Z(n13132) );
  COND1XL U11597 ( .A(n16939), .B(n12977), .C(n13132), .Z(n9937) );
  CANR2X1 U11598 ( .A(n12932), .B(poly14_shifted[279]), .C(n17655), .D(
        poly14_shifted[263]), .Z(n13133) );
  COND1XL U11599 ( .A(n16939), .B(n12932), .C(n13133), .Z(n10142) );
  CANR2X1 U11600 ( .A(n18018), .B(poly7_shifted[19]), .C(n17527), .D(
        Poly7[406]), .Z(n13134) );
  COND1XL U11601 ( .A(n16939), .B(n18018), .C(n13134), .Z(n10097) );
  CAN2X1 U11602 ( .A(n13189), .B(n13266), .Z(n13663) );
  CANR2X1 U11603 ( .A(n17750), .B(Poly8[71]), .C(n17620), .D(poly8_shifted[71]), .Z(n13135) );
  COND1XL U11604 ( .A(n16939), .B(n17750), .C(n13135), .Z(n11330) );
  CND2X1 U11605 ( .A(n12017), .B(n13136), .Z(n13137) );
  CANR2X1 U11606 ( .A(n17603), .B(poly13_shifted[358]), .C(n17640), .D(
        poly13_shifted[344]), .Z(n13138) );
  COND1XL U11607 ( .A(n16179), .B(n17603), .C(n13138), .Z(n10716) );
  CANR2X1 U11608 ( .A(n17603), .B(poly13_shifted[345]), .C(poly13_shifted[331]), .D(n16947), .Z(n13139) );
  COND1XL U11609 ( .A(n16605), .B(n17603), .C(n13139), .Z(n10729) );
  CENX1 U11610 ( .A(n14613), .B(n13140), .Z(n15187) );
  CEOXL U11611 ( .A(Poly4[58]), .B(Poly4[33]), .Z(n13141) );
  CENX1 U11612 ( .A(n15187), .B(n13141), .Z(n13143) );
  CMXI2XL U11613 ( .A0(n18210), .A1(Poly4[50]), .S(n12153), .Z(n13142) );
  COND1XL U11614 ( .A(n13143), .B(n15673), .C(n13142), .Z(n8806) );
  CANR2X1 U11615 ( .A(n12206), .B(poly7_shifted[371]), .C(n17449), .D(
        poly7_shifted[359]), .Z(n13144) );
  COND1XL U11616 ( .A(n16939), .B(n12206), .C(n13144), .Z(n9745) );
  CND2X1 U11617 ( .A(n13189), .B(n13145), .Z(n13146) );
  CANR2X1 U11618 ( .A(n17955), .B(poly9_shifted[83]), .C(n16702), .D(
        poly9_shifted[72]), .Z(n13147) );
  COND1XL U11619 ( .A(n17163), .B(n17955), .C(n13147), .Z(n11233) );
  CEOXL U11620 ( .A(Poly11[85]), .B(Poly11[31]), .Z(n13148) );
  CANR2X1 U11621 ( .A(n17683), .B(Poly11[46]), .C(n16919), .D(n13148), .Z(
        n13149) );
  COND1XL U11622 ( .A(n12764), .B(n17683), .C(n13149), .Z(n11143) );
  CIVX2 U11623 ( .A(n15673), .Z(n17598) );
  CANR2X1 U11624 ( .A(n18028), .B(poly7_shifted[307]), .C(n17598), .D(
        poly7_shifted[295]), .Z(n13150) );
  COND1XL U11625 ( .A(n16939), .B(n18028), .C(n13150), .Z(n9809) );
  CANR2X1 U11626 ( .A(n18028), .B(poly7_shifted[324]), .C(n17535), .D(
        poly7_shifted[312]), .Z(n13151) );
  COND1XL U11627 ( .A(n16179), .B(n18028), .C(n13151), .Z(n9792) );
  CIVX2 U11628 ( .A(n15673), .Z(n17453) );
  CANR2X1 U11629 ( .A(n12401), .B(poly7_shifted[403]), .C(n17453), .D(
        poly7_shifted[391]), .Z(n13152) );
  COND1XL U11630 ( .A(n17718), .B(n12401), .C(n13152), .Z(n9713) );
  CANR2X1 U11631 ( .A(n17217), .B(poly7_shifted[115]), .C(n17094), .D(
        poly7_shifted[103]), .Z(n13153) );
  COND1XL U11632 ( .A(n16939), .B(n17217), .C(n13153), .Z(n10001) );
  CND2X1 U11633 ( .A(n16700), .B(Poly6[51]), .Z(n14008) );
  CANR2X1 U11634 ( .A(n16063), .B(Poly6[50]), .C(Poly6[40]), .D(n14005), .Z(
        n13154) );
  COAN1X1 U11635 ( .A(n17567), .B(n14166), .C(n13154), .Z(n13155) );
  COND1XL U11636 ( .A(n14008), .B(Poly6[40]), .C(n13155), .Z(n9643) );
  CIVX2 U11637 ( .A(n15673), .Z(n16372) );
  CANR2X1 U11638 ( .A(n17053), .B(Poly1[199]), .C(n16372), .D(
        poly1_shifted[199]), .Z(n13156) );
  COND1XL U11639 ( .A(n16939), .B(n17053), .C(n13156), .Z(n9158) );
  COND1XL U11640 ( .A(poly3_shifted[15]), .B(n18206), .C(n18163), .Z(n13158)
         );
  CND2X1 U11641 ( .A(n15737), .B(poly3_shifted[29]), .Z(n13157) );
  COND1XL U11642 ( .A(n13158), .B(n15737), .C(n13157), .Z(n8925) );
  CIVX2 U11643 ( .A(n15648), .Z(n17449) );
  CANR2X1 U11644 ( .A(n18198), .B(poly1_shifted[314]), .C(n17449), .D(
        poly1_shifted[303]), .Z(n13159) );
  COND1XL U11645 ( .A(n17196), .B(n18198), .C(n13159), .Z(n9054) );
  CANR2X1 U11646 ( .A(n17574), .B(Poly7[238]), .C(n17705), .D(
        poly7_shifted[238]), .Z(n13160) );
  COND1XL U11647 ( .A(n12764), .B(n17574), .C(n13160), .Z(n9866) );
  CANR2X1 U11648 ( .A(n18018), .B(poly7_shifted[26]), .C(n17203), .D(
        poly7_shifted[14]), .Z(n13161) );
  COND1XL U11649 ( .A(n12764), .B(n18018), .C(n13161), .Z(n10090) );
  CANR2X1 U11650 ( .A(n17491), .B(poly13_shifted[522]), .C(n17634), .D(
        poly13_shifted[508]), .Z(n13162) );
  COND1XL U11651 ( .A(n11978), .B(n17491), .C(n13162), .Z(n10552) );
  CANR2X1 U11652 ( .A(n17491), .B(poly13_shifted[508]), .C(n17634), .D(
        poly13_shifted[494]), .Z(n13163) );
  COND1XL U11653 ( .A(n12764), .B(n17491), .C(n13163), .Z(n10566) );
  CND2X1 U11654 ( .A(n17755), .B(Poly10[41]), .Z(n16817) );
  CIVXL U11655 ( .A(Poly10[41]), .Z(n13164) );
  CANR11XL U11656 ( .A(n17317), .B(Poly10[25]), .C(n13164), .D(n11982), .Z(
        n13165) );
  COND1XL U11657 ( .A(Poly10[25]), .B(n16817), .C(n13165), .Z(n13166) );
  CMX2XL U11658 ( .A0(n13166), .A1(Poly10[37]), .S(n17411), .Z(n11066) );
  CANR2X1 U11659 ( .A(n18198), .B(poly1_shifted[327]), .C(n17613), .D(
        poly1_shifted[316]), .Z(n13167) );
  COND1XL U11660 ( .A(n11978), .B(n18198), .C(n13167), .Z(n9041) );
  CANR2X1 U11661 ( .A(n17332), .B(poly1_shifted[345]), .C(n18234), .D(
        poly1_shifted[334]), .Z(n13168) );
  COND1XL U11662 ( .A(n17699), .B(n17332), .C(n13168), .Z(n9023) );
  CANR2X1 U11663 ( .A(n17538), .B(poly0_shifted[156]), .C(Poly0[156]), .D(
        n17671), .Z(n13169) );
  COND1XL U11664 ( .A(n17674), .B(n11978), .C(n13169), .Z(n9421) );
  COND1XL U11665 ( .A(poly3_shifted[27]), .B(n18099), .C(n18098), .Z(n13171)
         );
  CND2X1 U11666 ( .A(n15737), .B(poly3_shifted[41]), .Z(n13170) );
  COND1XL U11667 ( .A(n13171), .B(n15737), .C(n13170), .Z(n8913) );
  CANR2X1 U11668 ( .A(n18028), .B(poly7_shifted[301]), .C(n17545), .D(
        poly7_shifted[289]), .Z(n13172) );
  COND1XL U11669 ( .A(n16950), .B(n18028), .C(n13172), .Z(n9815) );
  CANR2X1 U11670 ( .A(n17306), .B(Poly2[57]), .C(n17105), .D(poly2_shifted[57]), .Z(n13173) );
  COND1XL U11671 ( .A(n11997), .B(n17306), .C(n13173), .Z(n8953) );
  CANR2X1 U11672 ( .A(n12900), .B(poly13_shifted[52]), .C(n16427), .D(
        poly13_shifted[38]), .Z(n13174) );
  COND1XL U11673 ( .A(n17757), .B(n12900), .C(n13174), .Z(n11022) );
  CANR2X1 U11674 ( .A(n17603), .B(poly13_shifted[340]), .C(n17965), .D(
        poly13_shifted[326]), .Z(n13175) );
  COND1XL U11675 ( .A(n17757), .B(n17603), .C(n13175), .Z(n10734) );
  CANR2X1 U11676 ( .A(n17491), .B(poly13_shifted[500]), .C(n18234), .D(
        poly13_shifted[486]), .Z(n13176) );
  COND1XL U11677 ( .A(n16779), .B(n17491), .C(n13176), .Z(n10574) );
  CANR2X1 U11678 ( .A(n12210), .B(poly1_shifted[199]), .C(n16372), .D(
        poly1_shifted[188]), .Z(n13177) );
  COND1XL U11679 ( .A(n11978), .B(n12210), .C(n13177), .Z(n9169) );
  CANR2X1 U11680 ( .A(n17592), .B(poly13_shifted[276]), .C(n17634), .D(
        poly13_shifted[262]), .Z(n13178) );
  COND1XL U11681 ( .A(n16779), .B(n17592), .C(n13178), .Z(n10798) );
  CANR2X1 U11682 ( .A(n18028), .B(poly7_shifted[313]), .C(n17655), .D(
        poly7_shifted[301]), .Z(n13179) );
  COND1XL U11683 ( .A(n17090), .B(n18028), .C(n13179), .Z(n9803) );
  CANR2X1 U11684 ( .A(n18028), .B(poly7_shifted[311]), .C(n17285), .D(
        poly7_shifted[299]), .Z(n13180) );
  COND1XL U11685 ( .A(n16605), .B(n18028), .C(n13180), .Z(n9805) );
  CENX1 U11686 ( .A(dataselector[60]), .B(dataselector[7]), .Z(n13181) );
  CENX1 U11687 ( .A(n13181), .B(dataselector[63]), .Z(n13182) );
  CANR2X1 U11688 ( .A(n18160), .B(n17832), .C(n17280), .D(n13182), .Z(n13183)
         );
  COND1XL U11689 ( .A(n15799), .B(n15349), .C(n13183), .Z(n8781) );
  COND1XL U11690 ( .A(poly10_shifted[20]), .B(n18082), .C(n18200), .Z(n13184)
         );
  CMXI2XL U11691 ( .A0(n13185), .A1(n13184), .S(n13782), .Z(n11083) );
  CIVXL U11692 ( .A(Poly5[121]), .Z(n13187) );
  CANR2XL U11693 ( .A(n15574), .B(n18249), .C(poly5_shifted[121]), .D(n18017), 
        .Z(n13186) );
  COND1XL U11694 ( .A(n17031), .B(n13187), .C(n13186), .Z(n11405) );
  CANR2X1 U11695 ( .A(n17955), .B(poly9_shifted[86]), .C(n16702), .D(
        poly9_shifted[75]), .Z(n13188) );
  COND1XL U11696 ( .A(n16605), .B(n17955), .C(n13188), .Z(n11230) );
  CND2X1 U11697 ( .A(n13189), .B(n13227), .Z(n13190) );
  CNIVX8 U11698 ( .A(n13190), .Z(n17731) );
  CANR2X1 U11699 ( .A(n17731), .B(poly9_shifted[22]), .C(n18234), .D(
        poly9_shifted[11]), .Z(n13191) );
  COND1XL U11700 ( .A(n16605), .B(n17731), .C(n13191), .Z(n11294) );
  CANR2X1 U11701 ( .A(n12932), .B(poly14_shifted[283]), .C(n17174), .D(
        poly14_shifted[267]), .Z(n13192) );
  COND1XL U11702 ( .A(n16605), .B(n12932), .C(n13192), .Z(n10138) );
  CANR2X1 U11703 ( .A(n12211), .B(poly2_shifted[26]), .C(n17178), .D(
        poly2_shifted[14]), .Z(n13193) );
  COND1XL U11704 ( .A(n12764), .B(n12211), .C(n13193), .Z(n8996) );
  CANR2X1 U11705 ( .A(n13040), .B(poly7_shifted[343]), .C(n17453), .D(
        poly7_shifted[331]), .Z(n13194) );
  COND1XL U11706 ( .A(n16605), .B(n13040), .C(n13194), .Z(n9773) );
  CND2X1 U11707 ( .A(n17218), .B(n17826), .Z(n18153) );
  CIVX1 U11708 ( .A(n17076), .Z(n13522) );
  CANR2X1 U11709 ( .A(n17990), .B(poly13_shifted[479]), .C(poly13_shifted[465]), .D(n17755), .Z(n13195) );
  COND1XL U11710 ( .A(n17173), .B(n17990), .C(n13195), .Z(n10595) );
  CANR2X1 U11711 ( .A(n16842), .B(Poly4[54]), .C(n16840), .D(
        poly1_shifted[247]), .Z(n13199) );
  CANR2X1 U11712 ( .A(n16867), .B(Poly11[54]), .C(n16841), .D(
        poly1_shifted[275]), .Z(n13198) );
  CANR2X1 U11713 ( .A(n16877), .B(poly1_shifted[255]), .C(Poly6[28]), .D(
        n16837), .Z(n13197) );
  CANR2X1 U11714 ( .A(n16865), .B(poly5_shifted[36]), .C(n16861), .D(
        poly1_shifted[81]), .Z(n13196) );
  CAN4X1 U11715 ( .A(n13199), .B(n13198), .C(n13197), .D(n13196), .Z(n13216)
         );
  CANR2X1 U11716 ( .A(n16860), .B(poly13_shifted[365]), .C(n16843), .D(
        poly8_shifted[34]), .Z(n13203) );
  CANR2X1 U11717 ( .A(n16876), .B(poly7_shifted[230]), .C(n16838), .D(
        poly3_shifted[75]), .Z(n13202) );
  CANR2X1 U11718 ( .A(n16855), .B(poly0_shifted[68]), .C(n16853), .D(Poly6[27]), .Z(n13201) );
  CANR2X1 U11719 ( .A(n16863), .B(Poly3[49]), .C(n16852), .D(
        poly1_shifted[174]), .Z(n13200) );
  CAN4X1 U11720 ( .A(n13203), .B(n13202), .C(n13201), .D(n13200), .Z(n13215)
         );
  CANR2X1 U11721 ( .A(n16839), .B(poly3_shifted[74]), .C(n16862), .D(
        poly13_shifted[313]), .Z(n13207) );
  CANR2X1 U11722 ( .A(n12071), .B(poly10_shifted[42]), .C(Poly9[24]), .D(
        n16849), .Z(n13206) );
  CND2XL U11723 ( .A(n13493), .B(Poly6[48]), .Z(n13468) );
  CIVX2 U11724 ( .A(n13468), .Z(n13683) );
  CANR2X1 U11725 ( .A(n16844), .B(poly12_shifted[59]), .C(n13683), .D(n16873), 
        .Z(n13205) );
  CANR2X1 U11726 ( .A(n16864), .B(poly4_shifted[29]), .C(n16874), .D(
        Poly11[39]), .Z(n13204) );
  CAN4X1 U11727 ( .A(n13207), .B(n13206), .C(n13205), .D(n13204), .Z(n13214)
         );
  CNIVX4 U11728 ( .A(n13208), .Z(n16851) );
  CANR2X1 U11729 ( .A(n16875), .B(poly1_shifted[306]), .C(n16851), .D(
        poly7_shifted[52]), .Z(n13212) );
  CANR2X1 U11730 ( .A(n16850), .B(poly13_shifted[280]), .C(n16866), .D(
        poly7_shifted[380]), .Z(n13211) );
  CANR2X1 U11731 ( .A(n12084), .B(Poly2[60]), .C(n16872), .D(
        poly13_shifted[501]), .Z(n13210) );
  CANR2X1 U11732 ( .A(n12067), .B(poly7_shifted[379]), .C(n16854), .D(
        poly9_shifted[112]), .Z(n13209) );
  CAN4X1 U11733 ( .A(n13212), .B(n13211), .C(n13210), .D(n13209), .Z(n13213)
         );
  CND4X1 U11734 ( .A(n13216), .B(n13215), .C(n13214), .D(n13213), .Z(n13217)
         );
  CAOR2X2 U11735 ( .A(polydata[14]), .B(n17829), .C(n13217), .D(n16886), .Z(
        n8698) );
  CANR2X1 U11736 ( .A(n12192), .B(Poly1[233]), .C(n17527), .D(
        poly1_shifted[233]), .Z(n13218) );
  COND1XL U11737 ( .A(n17208), .B(n12192), .C(n13218), .Z(n9124) );
  CANR2X1 U11738 ( .A(n12192), .B(poly1_shifted[265]), .C(n17206), .D(
        poly1_shifted[254]), .Z(n13219) );
  COND1XL U11739 ( .A(n17004), .B(n12192), .C(n13219), .Z(n9103) );
  CANR2X1 U11740 ( .A(n12192), .B(poly1_shifted[262]), .C(n16435), .D(
        poly1_shifted[251]), .Z(n13220) );
  COND1XL U11741 ( .A(n17741), .B(n12192), .C(n13220), .Z(n9106) );
  CANR2X1 U11742 ( .A(n18018), .B(Poly7[20]), .C(n17266), .D(poly7_shifted[20]), .Z(n13221) );
  COND1XL U11743 ( .A(n17707), .B(n18018), .C(n13221), .Z(n10084) );
  CANR2X1 U11744 ( .A(n17053), .B(poly1_shifted[232]), .C(n17466), .D(
        poly1_shifted[221]), .Z(n13222) );
  COND1XL U11745 ( .A(n17185), .B(n17053), .C(n13222), .Z(n9136) );
  CIVX2 U11746 ( .A(n13223), .Z(n16801) );
  CIVXL U11747 ( .A(Poly1[228]), .Z(n13224) );
  CANR1XL U11748 ( .A(n16801), .B(n13224), .C(n18206), .Z(n13226) );
  CANR2X1 U11749 ( .A(n12192), .B(poly1_shifted[250]), .C(n13362), .D(
        Poly1[228]), .Z(n13225) );
  COND1XL U11750 ( .A(n13226), .B(n12192), .C(n13225), .Z(n9118) );
  CND2X4 U11751 ( .A(n12017), .B(n13227), .Z(n17615) );
  CANR2X1 U11752 ( .A(n17615), .B(poly13_shifted[333]), .C(n17755), .D(
        poly13_shifted[319]), .Z(n13228) );
  COND1XL U11753 ( .A(n17188), .B(n17615), .C(n13228), .Z(n10741) );
  CANR2X1 U11754 ( .A(n17987), .B(poly13_shifted[461]), .C(n17362), .D(
        poly13_shifted[447]), .Z(n13229) );
  COND1XL U11755 ( .A(n13482), .B(n17987), .C(n13229), .Z(n10613) );
  CANR2X1 U11756 ( .A(n13014), .B(poly13_shifted[202]), .C(n16919), .D(
        poly13_shifted[188]), .Z(n13230) );
  COND1XL U11757 ( .A(n11978), .B(n13014), .C(n13230), .Z(n10872) );
  CANR2X1 U11758 ( .A(n17603), .B(poly13_shifted[365]), .C(n17401), .D(
        poly13_shifted[351]), .Z(n13231) );
  COND1XL U11759 ( .A(n13482), .B(n17603), .C(n13231), .Z(n10709) );
  CANR2X1 U11760 ( .A(n17491), .B(poly13_shifted[525]), .C(poly13_shifted[511]), .D(n18017), .Z(n13232) );
  COND1XL U11761 ( .A(n13482), .B(n17491), .C(n13232), .Z(n10549) );
  COND1XL U11762 ( .A(poly13_shifted[313]), .B(n18249), .C(n18196), .Z(n13234)
         );
  CND2X1 U11763 ( .A(n17615), .B(poly13_shifted[327]), .Z(n13233) );
  COND1XL U11764 ( .A(n13234), .B(n17615), .C(n13233), .Z(n10747) );
  CANR2X1 U11765 ( .A(n17615), .B(poly13_shifted[330]), .C(n17640), .D(
        poly13_shifted[316]), .Z(n13235) );
  COND1XL U11766 ( .A(n11978), .B(n17615), .C(n13235), .Z(n10744) );
  CANR2X1 U11767 ( .A(n17615), .B(poly13_shifted[316]), .C(n17640), .D(
        poly13_shifted[302]), .Z(n13236) );
  COND1XL U11768 ( .A(n12764), .B(n17615), .C(n13236), .Z(n10758) );
  CANR2X1 U11769 ( .A(n12958), .B(poly14_shifted[80]), .C(n17655), .D(
        poly14_shifted[64]), .Z(n13237) );
  COND1XL U11770 ( .A(n12011), .B(n12958), .C(n13237), .Z(n10341) );
  CANR2X1 U11771 ( .A(n12287), .B(poly8_shifted[77]), .C(n18234), .D(
        poly8_shifted[63]), .Z(n13238) );
  COND1XL U11772 ( .A(n13482), .B(n12287), .C(n13238), .Z(n11338) );
  CND2X1 U11773 ( .A(n12017), .B(n13877), .Z(n13239) );
  CANR2X1 U11774 ( .A(n17969), .B(poly13_shifted[109]), .C(n17538), .D(
        poly13_shifted[95]), .Z(n13240) );
  COND1XL U11775 ( .A(n13482), .B(n17969), .C(n13240), .Z(n10965) );
  CIVX2 U11776 ( .A(n15673), .Z(n16488) );
  CANR2X1 U11777 ( .A(n17574), .B(poly7_shifted[237]), .C(n16488), .D(
        poly7_shifted[225]), .Z(n13241) );
  COND1XL U11778 ( .A(n16950), .B(n17574), .C(n13241), .Z(n9879) );
  CANR2X1 U11779 ( .A(n17977), .B(Poly13[158]), .C(n17755), .D(
        poly13_shifted[158]), .Z(n13242) );
  COND1XL U11780 ( .A(n17004), .B(n17977), .C(n13242), .Z(n10902) );
  CIVX2 U11781 ( .A(n18142), .Z(n17166) );
  CANR2X1 U11782 ( .A(n17574), .B(poly7_shifted[244]), .C(n16488), .D(
        poly7_shifted[232]), .Z(n13243) );
  COND1XL U11783 ( .A(n17166), .B(n17574), .C(n13243), .Z(n9872) );
  CANR2X1 U11784 ( .A(n13124), .B(poly13_shifted[31]), .C(n16479), .D(
        poly13_shifted[17]), .Z(n13244) );
  COND1XL U11785 ( .A(n17173), .B(n13124), .C(n13244), .Z(n11043) );
  CANR2X1 U11786 ( .A(n17977), .B(poly13_shifted[157]), .C(n17642), .D(
        poly13_shifted[143]), .Z(n13245) );
  COND1XL U11787 ( .A(n17196), .B(n17977), .C(n13245), .Z(n10917) );
  CIVXL U11788 ( .A(poly5_shifted[61]), .Z(n13247) );
  CANR2X1 U11789 ( .A(n12942), .B(n18206), .C(n17466), .D(poly5_shifted[47]), 
        .Z(n13246) );
  COND1XL U11790 ( .A(n17047), .B(n13247), .C(n13246), .Z(n11479) );
  CANR2X1 U11791 ( .A(n17047), .B(n13994), .C(n16488), .D(poly5_shifted[56]), 
        .Z(n13248) );
  COND1XL U11792 ( .A(n12942), .B(n13249), .C(n13248), .Z(n11470) );
  CANR2X1 U11793 ( .A(n17667), .B(poly13_shifted[237]), .C(n17504), .D(
        poly13_shifted[223]), .Z(n13250) );
  COND1XL U11794 ( .A(n13482), .B(n17667), .C(n13250), .Z(n10837) );
  CEOX1 U11795 ( .A(Poly3[77]), .B(Poly3[38]), .Z(n13252) );
  COAN1XL U11796 ( .A(n13252), .B(n13766), .C(n16391), .Z(n13254) );
  CANR2X1 U11797 ( .A(n17587), .B(Poly3[52]), .C(n13252), .D(n13251), .Z(
        n13253) );
  COND1XL U11798 ( .A(n13254), .B(n17262), .C(n13253), .Z(n8888) );
  CEOX1 U11799 ( .A(Poly3[49]), .B(Poly3[74]), .Z(n13256) );
  COAN1XL U11800 ( .A(n13256), .B(n16728), .C(n17188), .Z(n13258) );
  CANR2X1 U11801 ( .A(n17587), .B(poly3_shifted[77]), .C(n13256), .D(n13255), 
        .Z(n13257) );
  COND1XL U11802 ( .A(n13258), .B(n17262), .C(n13257), .Z(n8877) );
  CEOX1 U11803 ( .A(Poly3[73]), .B(Poly3[40]), .Z(n13259) );
  COAN1XL U11804 ( .A(n13259), .B(n13371), .C(n17753), .Z(n13261) );
  CAN2X1 U11805 ( .A(n18017), .B(n18208), .Z(n13372) );
  CANR2X1 U11806 ( .A(n17587), .B(Poly3[54]), .C(n13259), .D(n13372), .Z(
        n13260) );
  COND1XL U11807 ( .A(n13261), .B(n17262), .C(n13260), .Z(n8886) );
  CANR2X1 U11808 ( .A(n12192), .B(Poly1[228]), .C(n17094), .D(
        poly1_shifted[228]), .Z(n13262) );
  COND1XL U11809 ( .A(n12005), .B(n12192), .C(n13262), .Z(n9129) );
  CIVX2 U11810 ( .A(n12004), .Z(n17442) );
  CANR2X1 U11811 ( .A(n13124), .B(poly13_shifted[18]), .C(n17965), .D(
        Poly13[518]), .Z(n13263) );
  COND1XL U11812 ( .A(n17442), .B(n13124), .C(n13263), .Z(n11056) );
  CANR2X1 U11813 ( .A(n13014), .B(poly13_shifted[197]), .C(n17508), .D(
        poly13_shifted[183]), .Z(n13264) );
  COND1XL U11814 ( .A(n12000), .B(n13014), .C(n13264), .Z(n10877) );
  CANR2X1 U11815 ( .A(n14310), .B(Poly6[19]), .C(n17705), .D(poly6_shifted[19]), .Z(n13265) );
  COND1XL U11816 ( .A(n17658), .B(n14310), .C(n13265), .Z(n9674) );
  CANR2X1 U11817 ( .A(n12012), .B(poly1_shifted[90]), .C(n17705), .D(
        poly1_shifted[79]), .Z(n13268) );
  COND1XL U11818 ( .A(n17196), .B(n12012), .C(n13268), .Z(n9278) );
  CENX1 U11819 ( .A(Poly0[19]), .B(Poly0[216]), .Z(n13269) );
  COND1XL U11820 ( .A(n13269), .B(n17744), .C(n11985), .Z(n13271) );
  CMX2XL U11821 ( .A0(n13271), .A1(poly0_shifted[55]), .S(n13270), .Z(n9540)
         );
  CND2X1 U11822 ( .A(n12211), .B(poly2_shifted[17]), .Z(n13272) );
  COND4CXL U11823 ( .A(n17368), .B(n11993), .C(n12211), .D(n13272), .Z(n9005)
         );
  COND1XL U11824 ( .A(poly1_shifted[174]), .B(n18160), .C(n18159), .Z(n13274)
         );
  CND2X1 U11825 ( .A(n12210), .B(poly1_shifted[185]), .Z(n13273) );
  COND1XL U11826 ( .A(n13274), .B(n12210), .C(n13273), .Z(n9183) );
  CNR2X1 U11827 ( .A(n18053), .B(n16801), .Z(n18130) );
  CAOR1XL U11828 ( .A(Poly1[56]), .B(n13275), .C(n18130), .Z(n13277) );
  CANR2X1 U11829 ( .A(n12012), .B(poly1_shifted[78]), .C(Poly1[56]), .D(n13362), .Z(n13276) );
  COND1XL U11830 ( .A(n12012), .B(n13277), .C(n13276), .Z(n9290) );
  CANR2X1 U11831 ( .A(n12210), .B(poly1_shifted[198]), .C(n17705), .D(
        poly1_shifted[187]), .Z(n13278) );
  COND1XL U11832 ( .A(n17741), .B(n12210), .C(n13278), .Z(n9170) );
  CANR2X1 U11833 ( .A(n12210), .B(poly1_shifted[186]), .C(n16919), .D(
        poly1_shifted[175]), .Z(n13279) );
  COND1XL U11834 ( .A(n17196), .B(n12210), .C(n13279), .Z(n9182) );
  CANR2X1 U11835 ( .A(n12210), .B(Poly1[161]), .C(n17755), .D(
        poly1_shifted[161]), .Z(n13280) );
  COND1XL U11836 ( .A(n17697), .B(n12210), .C(n13280), .Z(n9196) );
  CANR2X1 U11837 ( .A(n17043), .B(Poly13[400]), .C(n17640), .D(
        poly13_shifted[400]), .Z(n13281) );
  COND1XL U11838 ( .A(n17062), .B(n17043), .C(n13281), .Z(n10660) );
  CANR2X1 U11839 ( .A(n17610), .B(poly1_shifted[149]), .C(n16985), .D(
        poly1_shifted[138]), .Z(n13282) );
  COND1XL U11840 ( .A(n12014), .B(n17610), .C(n13282), .Z(n9219) );
  COND1XL U11841 ( .A(n13522), .B(poly1_shifted[177]), .C(n18193), .Z(n13284)
         );
  CND2X1 U11842 ( .A(n12210), .B(poly1_shifted[188]), .Z(n13283) );
  COND1XL U11843 ( .A(n13284), .B(n12210), .C(n13283), .Z(n9180) );
  COND1XL U11844 ( .A(n13522), .B(poly1_shifted[81]), .C(n18193), .Z(n13286)
         );
  CND2X1 U11845 ( .A(n12012), .B(poly1_shifted[92]), .Z(n13285) );
  COND1XL U11846 ( .A(n13286), .B(n12012), .C(n13285), .Z(n9276) );
  CIVX2 U11847 ( .A(n15648), .Z(n17552) );
  CANR2X1 U11848 ( .A(n17043), .B(poly13_shifted[429]), .C(n17552), .D(
        poly13_shifted[415]), .Z(n13287) );
  COND1XL U11849 ( .A(n13482), .B(n17043), .C(n13287), .Z(n10645) );
  CANR2X1 U11850 ( .A(n12009), .B(poly14_shifted[129]), .C(n17508), .D(
        poly14_shifted[113]), .Z(n13288) );
  COND1XL U11851 ( .A(n17173), .B(n12009), .C(n13288), .Z(n10292) );
  CIVX2 U11852 ( .A(n15648), .Z(n16427) );
  CANR2X1 U11853 ( .A(n12009), .B(poly14_shifted[118]), .C(n16427), .D(
        poly14_shifted[102]), .Z(n13289) );
  COND1XL U11854 ( .A(n16779), .B(n12009), .C(n13289), .Z(n10303) );
  COND1XL U11855 ( .A(poly14_shifted[118]), .B(n18034), .C(n18088), .Z(n13291)
         );
  CND2X1 U11856 ( .A(n12009), .B(poly14_shifted[134]), .Z(n13290) );
  COND1XL U11857 ( .A(n13291), .B(n12009), .C(n13290), .Z(n10287) );
  CANR2X1 U11858 ( .A(n17610), .B(poly1_shifted[155]), .C(n16372), .D(
        poly1_shifted[144]), .Z(n13292) );
  COND1XL U11859 ( .A(n17062), .B(n17610), .C(n13292), .Z(n9213) );
  CEOXL U11860 ( .A(Poly8[86]), .B(Poly8[71]), .Z(n13293) );
  CANR2X1 U11861 ( .A(n17750), .B(Poly8[85]), .C(n17620), .D(n13293), .Z(
        n13294) );
  COND1XL U11862 ( .A(n17036), .B(n17750), .C(n13294), .Z(n11316) );
  CANR2X1 U11863 ( .A(n17750), .B(Poly8[79]), .C(n17121), .D(poly8_shifted[79]), .Z(n13295) );
  COND1XL U11864 ( .A(n17196), .B(n17750), .C(n13295), .Z(n11322) );
  CIVXL U11865 ( .A(Poly1[154]), .Z(n13296) );
  CANR1XL U11866 ( .A(n16801), .B(n13296), .C(n11996), .Z(n13298) );
  CANR2X1 U11867 ( .A(n12210), .B(poly1_shifted[176]), .C(n13362), .D(
        Poly1[154]), .Z(n13297) );
  COND1XL U11868 ( .A(n13298), .B(n12210), .C(n13297), .Z(n9192) );
  CENX1 U11869 ( .A(n14017), .B(n18239), .Z(n16380) );
  CENX1 U11870 ( .A(dataselector[62]), .B(dataselector[35]), .Z(n13299) );
  CENX1 U11871 ( .A(n16380), .B(n13299), .Z(n13302) );
  CND2XL U11872 ( .A(n16350), .B(dataselector[42]), .Z(n13301) );
  CND2XL U11873 ( .A(n12013), .B(n18248), .Z(n13300) );
  COND3XL U11874 ( .A(n13302), .B(n17959), .C(n13301), .D(n13300), .Z(n8753)
         );
  CANR2X1 U11875 ( .A(n13124), .B(poly13_shifted[45]), .C(n17238), .D(
        poly13_shifted[31]), .Z(n13303) );
  COND1XL U11876 ( .A(n13482), .B(n13124), .C(n13303), .Z(n11029) );
  CEOXL U11877 ( .A(n13796), .B(dataselector[52]), .Z(n13306) );
  CND2XL U11878 ( .A(n18099), .B(n18248), .Z(n13305) );
  CND2XL U11879 ( .A(dataselector[59]), .B(n16350), .Z(n13304) );
  COND3XL U11880 ( .A(n13306), .B(n17495), .C(n13305), .D(n13304), .Z(n8736)
         );
  CANR2XL U11881 ( .A(n12210), .B(poly1_shifted[193]), .C(n17206), .D(
        poly1_shifted[182]), .Z(n13307) );
  COND1XL U11882 ( .A(n17001), .B(n12210), .C(n13307), .Z(n9175) );
  CANR2X1 U11883 ( .A(n17043), .B(Poly13[396]), .C(n17545), .D(
        poly13_shifted[396]), .Z(n13308) );
  COND1XL U11884 ( .A(n17087), .B(n17043), .C(n13308), .Z(n10664) );
  CANR2X1 U11885 ( .A(n17043), .B(Poly13[392]), .C(n16427), .D(
        poly13_shifted[392]), .Z(n13309) );
  COND1XL U11886 ( .A(n17163), .B(n17043), .C(n13309), .Z(n10668) );
  CANR2X1 U11887 ( .A(n12210), .B(poly1_shifted[201]), .C(n17598), .D(
        poly1_shifted[190]), .Z(n13310) );
  COND1XL U11888 ( .A(n17004), .B(n12210), .C(n13310), .Z(n9167) );
  CIVX2 U11889 ( .A(n17259), .Z(n16583) );
  CEOXL U11890 ( .A(Poly13[524]), .B(Poly13[397]), .Z(n13311) );
  CANR2X1 U11891 ( .A(n17043), .B(poly13_shifted[425]), .C(n16583), .D(n13311), 
        .Z(n13312) );
  COND1XL U11892 ( .A(n17741), .B(n17043), .C(n13312), .Z(n10649) );
  CANR2X1 U11893 ( .A(n18198), .B(poly1_shifted[326]), .C(n17072), .D(
        poly1_shifted[315]), .Z(n13313) );
  COND1XL U11894 ( .A(n17741), .B(n18198), .C(n13313), .Z(n9042) );
  CANR2X1 U11895 ( .A(n18198), .B(poly1_shifted[328]), .C(n17620), .D(
        poly1_shifted[317]), .Z(n13314) );
  COND1XL U11896 ( .A(n17185), .B(n18198), .C(n13314), .Z(n9040) );
  CANR2X1 U11897 ( .A(n18198), .B(poly1_shifted[329]), .C(n17099), .D(
        poly1_shifted[318]), .Z(n13315) );
  COND1XL U11898 ( .A(n17004), .B(n18198), .C(n13315), .Z(n9039) );
  COND1XL U11899 ( .A(poly7_shifted[224]), .B(n12010), .C(n18185), .Z(n13317)
         );
  CND2XL U11900 ( .A(n17574), .B(poly7_shifted[236]), .Z(n13316) );
  COND1XL U11901 ( .A(n13317), .B(n17574), .C(n13316), .Z(n9880) );
  CIVX2 U11902 ( .A(n15648), .Z(n17466) );
  CANR2X1 U11903 ( .A(n17043), .B(Poly13[391]), .C(n17466), .D(
        poly13_shifted[391]), .Z(n13318) );
  COND1XL U11904 ( .A(n16939), .B(n17043), .C(n13318), .Z(n10669) );
  CANR2X1 U11905 ( .A(n16425), .B(poly1_shifted[124]), .C(n17705), .D(
        poly1_shifted[113]), .Z(n13319) );
  COND1XL U11906 ( .A(n17173), .B(n16425), .C(n13319), .Z(n9244) );
  CANR2XL U11907 ( .A(n16425), .B(poly1_shifted[132]), .C(n18017), .D(
        poly1_shifted[121]), .Z(n13320) );
  COND1XL U11908 ( .A(n17200), .B(n16425), .C(n13320), .Z(n9236) );
  COND1XL U11909 ( .A(poly14_shifted[133]), .B(n11986), .C(n18134), .Z(n13322)
         );
  CND2X1 U11910 ( .A(n12008), .B(poly14_shifted[149]), .Z(n13321) );
  COND1XL U11911 ( .A(n13322), .B(n12008), .C(n13321), .Z(n10272) );
  CANR2X1 U11912 ( .A(n17043), .B(Poly13[398]), .C(n16702), .D(
        poly13_shifted[398]), .Z(n13323) );
  COND1XL U11913 ( .A(n12764), .B(n17043), .C(n13323), .Z(n10662) );
  CANR2X1 U11914 ( .A(n12185), .B(Poly11[31]), .C(n17598), .D(
        poly11_shifted[31]), .Z(n13324) );
  COND1XL U11915 ( .A(n13482), .B(n12185), .C(n13324), .Z(n11158) );
  CENX1 U11916 ( .A(Poly4[44]), .B(n13329), .Z(n14615) );
  CEOX1 U11917 ( .A(n14615), .B(n15186), .Z(n13858) );
  CENX1 U11918 ( .A(Poly4[56]), .B(n18214), .Z(n16907) );
  CENX1 U11919 ( .A(Poly4[30]), .B(n16907), .Z(n13325) );
  CENX1 U11920 ( .A(n13858), .B(n13325), .Z(n13326) );
  CNR2XL U11921 ( .A(n13326), .B(n17826), .Z(n13327) );
  CANR1XL U11922 ( .A(Poly4[47]), .B(n12153), .C(n13327), .Z(n13328) );
  COND1XL U11923 ( .A(n17196), .B(n12153), .C(n13328), .Z(n8809) );
  CEOX1 U11924 ( .A(n13329), .B(n15186), .Z(n14485) );
  CENX1 U11925 ( .A(n14485), .B(n16907), .Z(n15822) );
  CEOX1 U11926 ( .A(n15822), .B(Poly4[18]), .Z(n13330) );
  CNR2X1 U11927 ( .A(n17495), .B(n13330), .Z(n13331) );
  CANR1XL U11928 ( .A(Poly4[35]), .B(n12153), .C(n13331), .Z(n13332) );
  COND1XL U11929 ( .A(n13275), .B(n12153), .C(n13332), .Z(n8821) );
  CANR2X1 U11930 ( .A(n12192), .B(Poly1[230]), .C(n17178), .D(
        poly1_shifted[230]), .Z(n13333) );
  COND1XL U11931 ( .A(n17757), .B(n12192), .C(n13333), .Z(n9127) );
  CANR2X1 U11932 ( .A(n12192), .B(Poly1[225]), .C(n17755), .D(
        poly1_shifted[225]), .Z(n13334) );
  COND1XL U11933 ( .A(n17697), .B(n12192), .C(n13334), .Z(n9132) );
  CANR2X1 U11934 ( .A(n18198), .B(poly1_shifted[305]), .C(n17215), .D(
        poly1_shifted[294]), .Z(n13335) );
  COND1XL U11935 ( .A(n16779), .B(n18198), .C(n13335), .Z(n9063) );
  CANR2X1 U11936 ( .A(n17610), .B(poly1_shifted[151]), .C(n17755), .D(
        poly1_shifted[140]), .Z(n13336) );
  COND1XL U11937 ( .A(n17087), .B(n17610), .C(n13336), .Z(n9217) );
  COND1XL U11938 ( .A(poly1_shifted[189]), .B(n18228), .C(n18227), .Z(n13338)
         );
  CND2X1 U11939 ( .A(n12210), .B(poly1_shifted[200]), .Z(n13337) );
  COND1XL U11940 ( .A(n13338), .B(n12210), .C(n13337), .Z(n9168) );
  CND2XL U11941 ( .A(n13275), .B(n17495), .Z(n18111) );
  COND1XL U11942 ( .A(poly1_shifted[131]), .B(n18053), .C(n18111), .Z(n13340)
         );
  CND2X1 U11943 ( .A(n17610), .B(poly1_shifted[142]), .Z(n13339) );
  COND1XL U11944 ( .A(n13340), .B(n17610), .C(n13339), .Z(n9226) );
  CANR2X1 U11945 ( .A(n12210), .B(poly1_shifted[192]), .C(n16644), .D(
        poly1_shifted[181]), .Z(n13341) );
  COND1XL U11946 ( .A(n12006), .B(n12210), .C(n13341), .Z(n9176) );
  CANR2X1 U11947 ( .A(n17610), .B(Poly1[156]), .C(n17705), .D(
        poly1_shifted[156]), .Z(n13342) );
  COND1XL U11948 ( .A(n11978), .B(n17610), .C(n13342), .Z(n9201) );
  CND2X1 U11949 ( .A(n17935), .B(poly5_shifted[69]), .Z(n13344) );
  CND2XL U11950 ( .A(n17965), .B(poly5_shifted[55]), .Z(n13343) );
  COND3XL U11951 ( .A(n15378), .B(n12000), .C(n13344), .D(n13343), .Z(n11471)
         );
  CIVXL U11952 ( .A(Poly12[89]), .Z(n13345) );
  CANR1XL U11953 ( .A(n17994), .B(n13345), .C(n18189), .Z(n13347) );
  CIVX4 U11954 ( .A(n18001), .Z(n17652) );
  CANR2X1 U11955 ( .A(n17652), .B(poly12_shifted[121]), .C(n17995), .D(
        Poly12[89]), .Z(n13346) );
  COND1XL U11956 ( .A(n13347), .B(n17652), .C(n13346), .Z(n10427) );
  CANR2X1 U11957 ( .A(n12299), .B(poly1_shifted[59]), .C(n17063), .D(
        poly1_shifted[48]), .Z(n13348) );
  COND1XL U11958 ( .A(n17062), .B(n12299), .C(n13348), .Z(n9309) );
  CANR2X1 U11959 ( .A(n12299), .B(Poly1[61]), .C(n18234), .D(poly1_shifted[61]), .Z(n13349) );
  COND1XL U11960 ( .A(n17185), .B(n12299), .C(n13349), .Z(n9296) );
  CANR2X1 U11961 ( .A(n12299), .B(Poly1[59]), .C(n18234), .D(poly1_shifted[59]), .Z(n13350) );
  COND1XL U11962 ( .A(n17741), .B(n12299), .C(n13350), .Z(n9298) );
  CANR2X1 U11963 ( .A(n13351), .B(poly9_shifted[74]), .C(n17560), .D(
        poly9_shifted[63]), .Z(n13352) );
  COND1XL U11964 ( .A(n13482), .B(n13351), .C(n13352), .Z(n11242) );
  CANR2X1 U11965 ( .A(n18198), .B(poly1_shifted[315]), .C(n17705), .D(
        poly1_shifted[304]), .Z(n13353) );
  COND1XL U11966 ( .A(n17211), .B(n18198), .C(n13353), .Z(n9053) );
  CIVX2 U11967 ( .A(n15648), .Z(n17401) );
  CANR2X1 U11968 ( .A(n17043), .B(Poly13[393]), .C(n17401), .D(
        poly13_shifted[393]), .Z(n13355) );
  COND1XL U11969 ( .A(n17208), .B(n17043), .C(n13355), .Z(n10667) );
  CEOXL U11970 ( .A(Poly13[527]), .B(Poly13[400]), .Z(n13356) );
  CANR2X1 U11971 ( .A(n17043), .B(poly13_shifted[428]), .C(n16787), .D(n13356), 
        .Z(n13357) );
  COND1XL U11972 ( .A(n17004), .B(n17043), .C(n13357), .Z(n10646) );
  CANR2X1 U11973 ( .A(n17043), .B(Poly13[397]), .C(n17508), .D(
        poly13_shifted[397]), .Z(n13358) );
  COND1XL U11974 ( .A(n17065), .B(n17043), .C(n13358), .Z(n10663) );
  CANR2X1 U11975 ( .A(n17043), .B(poly13_shifted[399]), .C(poly13_shifted[385]), .D(n18017), .Z(n13359) );
  COND1XL U11976 ( .A(n17697), .B(n17043), .C(n13359), .Z(n10675) );
  CANR2X1 U11977 ( .A(n17750), .B(poly8_shifted[80]), .C(n17545), .D(
        poly8_shifted[66]), .Z(n13360) );
  COND1XL U11978 ( .A(n16775), .B(n17750), .C(n13360), .Z(n11335) );
  CIVXL U11979 ( .A(Poly1[201]), .Z(n13361) );
  CANR1XL U11980 ( .A(n16801), .B(n13361), .C(n18082), .Z(n13364) );
  CANR2X1 U11981 ( .A(n17053), .B(poly1_shifted[223]), .C(n13362), .D(
        Poly1[201]), .Z(n13363) );
  COND1XL U11982 ( .A(n13364), .B(n17053), .C(n13363), .Z(n9145) );
  CANR2X1 U11983 ( .A(n17610), .B(Poly1[154]), .C(n17504), .D(
        poly1_shifted[154]), .Z(n13365) );
  COND1XL U11984 ( .A(n17305), .B(n17610), .C(n13365), .Z(n9203) );
  CANR2X1 U11985 ( .A(n18198), .B(poly1_shifted[325]), .C(n17449), .D(
        poly1_shifted[314]), .Z(n13366) );
  COND1XL U11986 ( .A(n17305), .B(n18198), .C(n13366), .Z(n9043) );
  CANR2X1 U11987 ( .A(n12192), .B(poly1_shifted[261]), .C(n17063), .D(
        poly1_shifted[250]), .Z(n13368) );
  COND1XL U11988 ( .A(n17735), .B(n12192), .C(n13368), .Z(n9107) );
  COND1XL U11989 ( .A(poly1_shifted[247]), .B(n11999), .C(n18203), .Z(n13370)
         );
  CND2X1 U11990 ( .A(n12192), .B(poly1_shifted[258]), .Z(n13369) );
  COND1XL U11991 ( .A(n13370), .B(n12192), .C(n13369), .Z(n9110) );
  COAN1XL U11992 ( .A(Poly3[54]), .B(n13371), .C(n12005), .Z(n13374) );
  CANR2X1 U11993 ( .A(n13372), .B(Poly3[54]), .C(n17359), .D(poly3_shifted[82]), .Z(n13373) );
  COND1XL U11994 ( .A(n17359), .B(n13374), .C(n13373), .Z(n8872) );
  CAN2XL U11995 ( .A(n18017), .B(poly1_shifted[55]), .Z(n13375) );
  CANR1XL U11996 ( .A(Poly1[55]), .B(n12299), .C(n13375), .Z(n13376) );
  COND1XL U11997 ( .A(n12296), .B(n12299), .C(n13376), .Z(n9302) );
  CENX2 U11998 ( .A(Poly4[57]), .B(n14614), .Z(n16068) );
  CENX1 U11999 ( .A(n13800), .B(n16068), .Z(n16988) );
  CENX1 U12000 ( .A(Poly4[20]), .B(n16988), .Z(n13377) );
  CNR2XL U12001 ( .A(n17744), .B(n13377), .Z(n13378) );
  CANR1XL U12002 ( .A(Poly4[37]), .B(n12153), .C(n13378), .Z(n13379) );
  COND1XL U12003 ( .A(n11987), .B(n12153), .C(n13379), .Z(n8819) );
  CANR2X1 U12004 ( .A(n18198), .B(poly1_shifted[303]), .C(n17449), .D(
        poly1_shifted[292]), .Z(n13380) );
  COND1XL U12005 ( .A(n17442), .B(n18198), .C(n13380), .Z(n9065) );
  CANR2X1 U12006 ( .A(n17332), .B(poly1_shifted[335]), .C(n16326), .D(
        poly1_shifted[324]), .Z(n13381) );
  COND1XL U12007 ( .A(n17417), .B(n17332), .C(n13381), .Z(n9033) );
  CANR2X1 U12008 ( .A(n17043), .B(Poly13[388]), .C(n16702), .D(
        poly13_shifted[388]), .Z(n13382) );
  COND1XL U12009 ( .A(n17423), .B(n17043), .C(n13382), .Z(n10672) );
  CANR2X1 U12010 ( .A(n12210), .B(poly1_shifted[194]), .C(n16787), .D(
        poly1_shifted[183]), .Z(n13383) );
  COND1XL U12011 ( .A(n12296), .B(n12210), .C(n13383), .Z(n9174) );
  CIVX2 U12012 ( .A(n18210), .Z(n17567) );
  CANR2X1 U12013 ( .A(n18198), .B(poly1_shifted[317]), .C(n17266), .D(
        poly1_shifted[306]), .Z(n13384) );
  COND1XL U12014 ( .A(n17567), .B(n18198), .C(n13384), .Z(n9051) );
  CANR2X1 U12015 ( .A(n12299), .B(poly1_shifted[61]), .C(n18234), .D(
        poly1_shifted[50]), .Z(n13385) );
  COND1XL U12016 ( .A(n17567), .B(n12299), .C(n13385), .Z(n9307) );
  CANR2X1 U12017 ( .A(n18198), .B(poly1_shifted[318]), .C(n17508), .D(
        poly1_shifted[307]), .Z(n13386) );
  COND1XL U12018 ( .A(n17664), .B(n18198), .C(n13386), .Z(n9050) );
  CIVX2 U12019 ( .A(n18176), .Z(n17673) );
  CANR2X1 U12020 ( .A(n17332), .B(Poly1[339]), .C(n17560), .D(
        poly1_shifted[339]), .Z(n13387) );
  COND1XL U12021 ( .A(n17673), .B(n17332), .C(n13387), .Z(n9018) );
  CEOXL U12022 ( .A(Poly13[516]), .B(Poly13[389]), .Z(n13388) );
  CANR2X1 U12023 ( .A(n17043), .B(poly13_shifted[417]), .C(n17105), .D(n13388), 
        .Z(n13389) );
  COND1XL U12024 ( .A(n17658), .B(n17043), .C(n13389), .Z(n10657) );
  CNIVX1 U12025 ( .A(n18257), .Z(n18324) );
  CNIVX1 U12026 ( .A(n18257), .Z(n18314) );
  CNIVX1 U12027 ( .A(n18257), .Z(n18291) );
  CNIVX1 U12028 ( .A(n18257), .Z(n18308) );
  CNIVX1 U12029 ( .A(n18257), .Z(n18317) );
  CNIVX1 U12030 ( .A(n18257), .Z(n18306) );
  CNIVX1 U12031 ( .A(n18257), .Z(n18372) );
  CNIVX1 U12032 ( .A(n18257), .Z(n18325) );
  CNIVX1 U12033 ( .A(n18257), .Z(n18336) );
  CNIVX1 U12034 ( .A(n18257), .Z(n18318) );
  CNIVX1 U12035 ( .A(n18257), .Z(n18333) );
  CNIVX1 U12036 ( .A(n18257), .Z(n18337) );
  CNIVX1 U12037 ( .A(n18257), .Z(n18361) );
  CNIVX1 U12038 ( .A(n18257), .Z(n18330) );
  CNIVX1 U12039 ( .A(n18257), .Z(n18265) );
  CNIVX1 U12040 ( .A(n18257), .Z(n18264) );
  CNIVX1 U12041 ( .A(n18257), .Z(n18299) );
  CNIVX1 U12042 ( .A(n18257), .Z(n18373) );
  CNIVX1 U12043 ( .A(n18257), .Z(n18393) );
  CNIVX1 U12044 ( .A(n18257), .Z(n18358) );
  CNIVX1 U12045 ( .A(n18257), .Z(n18322) );
  CNIVX1 U12046 ( .A(n18257), .Z(n18328) );
  CNIVX1 U12047 ( .A(n18257), .Z(n18339) );
  CNIVX1 U12048 ( .A(n18257), .Z(n18349) );
  CNIVX1 U12049 ( .A(n18257), .Z(n18394) );
  CNIVX1 U12050 ( .A(n18257), .Z(n18395) );
  CNIVX1 U12051 ( .A(n18257), .Z(n18298) );
  CNIVX1 U12052 ( .A(n18257), .Z(n18263) );
  CNIVX1 U12053 ( .A(n18257), .Z(n18259) );
  CNIVX1 U12054 ( .A(n18257), .Z(n18355) );
  CNIVX1 U12055 ( .A(n18257), .Z(n18320) );
  CNIVX1 U12056 ( .A(n18257), .Z(n18357) );
  CNIVX1 U12057 ( .A(n18257), .Z(n18296) );
  CNIVX1 U12058 ( .A(n18257), .Z(n18362) );
  CNIVX1 U12059 ( .A(n18257), .Z(n18363) );
  CNIVX1 U12060 ( .A(n18257), .Z(n18364) );
  CNIVX1 U12061 ( .A(n18257), .Z(n18365) );
  CNIVX1 U12062 ( .A(n18257), .Z(n18295) );
  CNIVX1 U12063 ( .A(n18257), .Z(n18366) );
  CNIVX1 U12064 ( .A(n18257), .Z(n18367) );
  CNIVX1 U12065 ( .A(n18257), .Z(n18287) );
  CNIVX1 U12066 ( .A(n18257), .Z(n18374) );
  CNIVX1 U12067 ( .A(n18257), .Z(n18375) );
  CNIVX1 U12068 ( .A(n18257), .Z(n18274) );
  CNIVX1 U12069 ( .A(n18257), .Z(n18376) );
  CNIVX1 U12070 ( .A(n18257), .Z(n18382) );
  CNIVX1 U12071 ( .A(n18257), .Z(n18275) );
  CNIVX1 U12072 ( .A(n18257), .Z(n18277) );
  CNIVX1 U12073 ( .A(n18257), .Z(n18356) );
  CNIVX1 U12074 ( .A(n18257), .Z(n18278) );
  CNIVX1 U12075 ( .A(n18257), .Z(n18283) );
  CNIVX1 U12076 ( .A(n18257), .Z(n18302) );
  CNIVX1 U12077 ( .A(n18257), .Z(n18344) );
  CNIVX1 U12078 ( .A(n18257), .Z(n18288) );
  CNIVX1 U12079 ( .A(n18257), .Z(n18369) );
  CNIVX1 U12080 ( .A(n18257), .Z(n18270) );
  CNIVX1 U12081 ( .A(n18257), .Z(n18340) );
  CNIVX1 U12082 ( .A(n18257), .Z(n18286) );
  CNIVX1 U12083 ( .A(n18257), .Z(n18290) );
  CNIVX1 U12084 ( .A(n18257), .Z(n18293) );
  CNIVX1 U12085 ( .A(n18257), .Z(n18399) );
  CNIVX1 U12086 ( .A(n18257), .Z(n18294) );
  CNIVX1 U12087 ( .A(n18257), .Z(n18297) );
  CNIVX1 U12088 ( .A(n18257), .Z(n18303) );
  CNIVX1 U12089 ( .A(n18257), .Z(n18304) );
  CNIVX1 U12090 ( .A(n18257), .Z(n18307) );
  CNIVX1 U12091 ( .A(n18257), .Z(n18309) );
  CNIVX1 U12092 ( .A(n18257), .Z(n18313) );
  CNIVX1 U12093 ( .A(n18257), .Z(n18377) );
  CNIVX1 U12094 ( .A(n18257), .Z(n18319) );
  CNIVX1 U12095 ( .A(n18257), .Z(n18321) );
  CNIVX1 U12096 ( .A(n18257), .Z(n18385) );
  CNIVX1 U12097 ( .A(n18257), .Z(n18326) );
  CNIVX1 U12098 ( .A(n18257), .Z(n18327) );
  CNIVX1 U12099 ( .A(n18257), .Z(n18329) );
  CNIVX1 U12100 ( .A(n18257), .Z(n18331) );
  CNIVX1 U12101 ( .A(n18257), .Z(n18332) );
  CNIVX1 U12102 ( .A(n18257), .Z(n18315) );
  CNIVX1 U12103 ( .A(n18257), .Z(n18334) );
  CNIVX1 U12104 ( .A(n18257), .Z(n18401) );
  CNIVX1 U12105 ( .A(n18257), .Z(n18335) );
  CNIVX1 U12106 ( .A(n18257), .Z(n18397) );
  CNIVX1 U12107 ( .A(n18257), .Z(n18338) );
  CNIVX1 U12108 ( .A(n18257), .Z(n18396) );
  CNIVX1 U12109 ( .A(n18257), .Z(n18387) );
  CNIVX1 U12110 ( .A(n18257), .Z(n18388) );
  CNIVX1 U12111 ( .A(n18257), .Z(n18351) );
  CNIVX1 U12112 ( .A(n18257), .Z(n18386) );
  CNIVX1 U12113 ( .A(n18257), .Z(n18352) );
  CNIVX1 U12114 ( .A(n18257), .Z(n18353) );
  CNIVX1 U12115 ( .A(n18257), .Z(n18289) );
  CNIVX1 U12116 ( .A(n18257), .Z(n18323) );
  CNIVX1 U12117 ( .A(n18257), .Z(n18343) );
  CNIVX1 U12118 ( .A(n18257), .Z(n18342) );
  CNIVX1 U12119 ( .A(n18257), .Z(n18370) );
  CNIVX1 U12120 ( .A(n18257), .Z(n18371) );
  CNIVX1 U12121 ( .A(n18257), .Z(n18383) );
  CNIVX1 U12122 ( .A(n18257), .Z(n18380) );
  CNIVX1 U12123 ( .A(n18257), .Z(n18262) );
  CNIVX1 U12124 ( .A(n18257), .Z(n18292) );
  CNIVX1 U12125 ( .A(n18257), .Z(n18276) );
  CNIVX1 U12126 ( .A(n18257), .Z(n18316) );
  CNIVX1 U12127 ( .A(n18257), .Z(n18368) );
  CNIVX1 U12128 ( .A(n18257), .Z(n18359) );
  CNIVX1 U12129 ( .A(n18257), .Z(n18384) );
  CNIVX1 U12130 ( .A(n18257), .Z(n18398) );
  CNIVX1 U12131 ( .A(n18257), .Z(n18305) );
  CNIVX1 U12132 ( .A(n18257), .Z(n18381) );
  CNIVX1 U12133 ( .A(n18257), .Z(n18390) );
  CNIVX1 U12134 ( .A(n18257), .Z(n18402) );
  CNIVX1 U12135 ( .A(n18257), .Z(n18341) );
  CNIVX1 U12136 ( .A(n18257), .Z(n18379) );
  CNIVX1 U12137 ( .A(n18257), .Z(n18266) );
  CNIVX1 U12138 ( .A(n18257), .Z(n18350) );
  CNIVX1 U12139 ( .A(n18257), .Z(n18267) );
  CNIVX1 U12140 ( .A(n18257), .Z(n18312) );
  CNIVX1 U12141 ( .A(n18257), .Z(n18311) );
  CNIVX1 U12142 ( .A(n18257), .Z(n18268) );
  CNIVX1 U12143 ( .A(n18257), .Z(n18281) );
  CNIVX1 U12144 ( .A(n18257), .Z(n18269) );
  CNIVX1 U12145 ( .A(n18257), .Z(n18391) );
  CNIVX1 U12146 ( .A(n18257), .Z(n18258) );
  CNIVX1 U12147 ( .A(n18257), .Z(n18360) );
  CNIVX1 U12148 ( .A(n18257), .Z(n18300) );
  CNIVX1 U12149 ( .A(n18257), .Z(n18271) );
  CNIVX1 U12150 ( .A(n18257), .Z(n18310) );
  CNIVX1 U12151 ( .A(n18257), .Z(n18284) );
  CNIVX1 U12152 ( .A(n18257), .Z(n18261) );
  CNIVX1 U12153 ( .A(n18257), .Z(n18301) );
  CNIVX1 U12154 ( .A(n18257), .Z(n18260) );
  CNIVX1 U12155 ( .A(n18257), .Z(n18389) );
  CNIVX1 U12156 ( .A(n18257), .Z(n18272) );
  CNIVX1 U12157 ( .A(n18257), .Z(n18392) );
  CNIVX1 U12158 ( .A(n18257), .Z(n18378) );
  CNIVX1 U12159 ( .A(n18257), .Z(n18280) );
  CNIVX1 U12160 ( .A(n18257), .Z(n18346) );
  CNIVX1 U12161 ( .A(n18257), .Z(n18273) );
  CNIVX1 U12162 ( .A(n18257), .Z(n18400) );
  CNIVX1 U12163 ( .A(n18257), .Z(n18282) );
  CNIVX1 U12164 ( .A(n18257), .Z(n18348) );
  CNIVX1 U12165 ( .A(n18257), .Z(n18345) );
  CNIVX1 U12166 ( .A(n18257), .Z(n18279) );
  CNIVX1 U12167 ( .A(n18257), .Z(n18285) );
  CNIVX1 U12168 ( .A(n18257), .Z(n18354) );
  CNIVX1 U12169 ( .A(n18257), .Z(n18347) );
  CMXI2X1 U12170 ( .A0(n18189), .A1(poly12_shifted[25]), .S(n12997), .Z(n13390) );
  CND2X1 U12171 ( .A(n17755), .B(Poly12[120]), .Z(n14287) );
  CND2X1 U12172 ( .A(n13390), .B(n14287), .Z(n10523) );
  CMXI2X1 U12173 ( .A0(n13428), .A1(poly12_shifted[18]), .S(n12997), .Z(n13391) );
  CND2X1 U12174 ( .A(n17755), .B(Poly12[113]), .Z(n14295) );
  CND2X1 U12175 ( .A(n13391), .B(n14295), .Z(n10530) );
  CEOXL U12176 ( .A(scrambler[24]), .B(scrambler[19]), .Z(n13392) );
  CENX1 U12177 ( .A(n17882), .B(n13392), .Z(n17862) );
  CEOX1 U12178 ( .A(scrambler[18]), .B(scrambler[16]), .Z(n17868) );
  CENX1 U12179 ( .A(n17868), .B(scrambler[10]), .Z(n13393) );
  CENX1 U12180 ( .A(n17862), .B(n13393), .Z(dataout[26]) );
  CENX1 U12181 ( .A(Poly11[81]), .B(n15844), .Z(n13612) );
  COND1XL U12182 ( .A(Poly11[42]), .B(n13612), .C(n18017), .Z(n13395) );
  CIVDX2 U12183 ( .A(n17123), .Z0(n18249), .Z1(n17200) );
  CMXI2X1 U12184 ( .A0(n18249), .A1(Poly11[57]), .S(n17683), .Z(n13394) );
  COND4CX1 U12185 ( .A(n13612), .B(Poly11[42]), .C(n13395), .D(n13394), .Z(
        n11132) );
  CND2X1 U12186 ( .A(n17755), .B(Poly11[78]), .Z(n14303) );
  CND2X1 U12187 ( .A(n14300), .B(Poly11[48]), .Z(n13397) );
  CMXI2X1 U12188 ( .A0(n14436), .A1(Poly11[63]), .S(n17683), .Z(n13396) );
  COND3X1 U12189 ( .A(Poly11[48]), .B(n14303), .C(n13397), .D(n13396), .Z(
        n11126) );
  COND1XL U12190 ( .A(Poly9[108]), .B(Poly9[87]), .C(n17620), .Z(n13399) );
  CMXI2X1 U12191 ( .A0(n12415), .A1(poly9_shifted[109]), .S(n12262), .Z(n13398) );
  COND4CX1 U12192 ( .A(Poly9[87]), .B(Poly9[108]), .C(n13399), .D(n13398), .Z(
        n11207) );
  COND1XL U12193 ( .A(Poly9[106]), .B(Poly9[85]), .C(n17705), .Z(n13401) );
  CMXI2X1 U12194 ( .A0(n18108), .A1(poly9_shifted[107]), .S(n12262), .Z(n13400) );
  COND4CX1 U12195 ( .A(Poly9[85]), .B(Poly9[106]), .C(n13401), .D(n13400), .Z(
        n11209) );
  COND1XL U12196 ( .A(Poly9[109]), .B(Poly9[88]), .C(n17965), .Z(n13403) );
  CMXI2X1 U12197 ( .A0(n18053), .A1(poly9_shifted[110]), .S(n12262), .Z(n13402) );
  COND4CX1 U12198 ( .A(Poly9[88]), .B(Poly9[109]), .C(n13403), .D(n13402), .Z(
        n11206) );
  COND1XL U12199 ( .A(Poly12[111]), .B(Poly12[15]), .C(n17538), .Z(n13405) );
  CMXI2X1 U12200 ( .A0(n14436), .A1(Poly12[31]), .S(n12997), .Z(n13404) );
  COND4CX1 U12201 ( .A(Poly12[15]), .B(Poly12[111]), .C(n13405), .D(n13404), 
        .Z(n10501) );
  CENX1 U12202 ( .A(Poly11[82]), .B(n17680), .Z(n13563) );
  COND1XL U12203 ( .A(Poly11[43]), .B(n13563), .C(n17714), .Z(n13407) );
  CMXI2X1 U12204 ( .A0(n18095), .A1(Poly11[58]), .S(n17683), .Z(n13406) );
  COND4CX1 U12205 ( .A(n13563), .B(Poly11[43]), .C(n13407), .D(n13406), .Z(
        n11131) );
  CIVDX1 U12206 ( .A(n13481), .Z0(n13499), .Z1(n13408) );
  CND2X1 U12207 ( .A(n17932), .B(Poly5[2]), .Z(n13409) );
  COND4CX1 U12208 ( .A(n13410), .B(n16303), .C(n17932), .D(n13409), .Z(n11524)
         );
  COND1XL U12209 ( .A(poly2_shifted[16]), .B(n18167), .C(n18166), .Z(n13411)
         );
  CIVX1 U12210 ( .A(poly2_shifted[28]), .Z(n13434) );
  CMXI2X1 U12211 ( .A0(n13411), .A1(n13434), .S(n12211), .Z(n8994) );
  CMXI2X1 U12212 ( .A0(n13499), .A1(n13498), .S(Poly6[39]), .Z(n13413) );
  CMXI2X1 U12213 ( .A0(n14297), .A1(Poly6[49]), .S(n16063), .Z(n13412) );
  CND2X1 U12214 ( .A(n13413), .B(n13412), .Z(n9644) );
  CMXI2X1 U12215 ( .A0(n12010), .A1(Poly6[32]), .S(n16063), .Z(n13415) );
  CMXI2X1 U12216 ( .A0(n13499), .A1(n13498), .S(Poly6[22]), .Z(n13414) );
  CND2X1 U12217 ( .A(n13415), .B(n13414), .Z(n9661) );
  CND2X1 U12218 ( .A(n17932), .B(Poly5[1]), .Z(n13416) );
  COND4CX1 U12219 ( .A(n13417), .B(n17697), .C(n17932), .D(n13416), .Z(n11525)
         );
  CND2X1 U12220 ( .A(n17640), .B(Poly15[46]), .Z(n18040) );
  CIVDX1 U12221 ( .A(n13418), .Z0(n18105), .Z1(n17004) );
  COND4CXL U12222 ( .A(Poly11[39]), .B(n14300), .C(n18034), .D(n11998), .Z(
        n13423) );
  CND2X1 U12223 ( .A(n17747), .B(Poly11[54]), .Z(n13422) );
  COND3X1 U12224 ( .A(Poly11[39]), .B(n14303), .C(n13423), .D(n13422), .Z(
        n11135) );
  CND2X1 U12225 ( .A(n17930), .B(poly5_shifted[44]), .Z(n13425) );
  CND2X1 U12226 ( .A(n18234), .B(poly5_shifted[30]), .Z(n13424) );
  COND3X1 U12227 ( .A(n17932), .B(n17004), .C(n13425), .D(n13424), .Z(n11496)
         );
  CND2X1 U12228 ( .A(n17930), .B(poly5_shifted[43]), .Z(n13427) );
  CND2X1 U12229 ( .A(n17285), .B(poly5_shifted[29]), .Z(n13426) );
  COND3X1 U12230 ( .A(n17932), .B(n17185), .C(n13427), .D(n13426), .Z(n11497)
         );
  CNR2X1 U12231 ( .A(n13428), .B(n13683), .Z(n13429) );
  CIVX1 U12232 ( .A(Poly6[2]), .Z(n13686) );
  CMXI2X1 U12233 ( .A0(n13429), .A1(n13686), .S(n14310), .Z(n9691) );
  CND2XL U12234 ( .A(n11978), .B(n11972), .Z(n13430) );
  CMXI2XL U12235 ( .A0(dataselector[28]), .A1(n13430), .S(n17831), .Z(n13432)
         );
  CENX1 U12236 ( .A(n17830), .B(n14017), .Z(n18233) );
  CNR2XL U12237 ( .A(n18233), .B(n17495), .Z(n13431) );
  CMXI2X1 U12238 ( .A0(n13432), .A1(dataselector[21]), .S(n13431), .Z(n8767)
         );
  CND2X1 U12239 ( .A(n16999), .B(Poly2[65]), .Z(n14772) );
  CND2X1 U12240 ( .A(n12211), .B(poly2_shifted[19]), .Z(n13433) );
  COND4CX1 U12241 ( .A(n14772), .B(n17718), .C(n12211), .D(n13433), .Z(n9003)
         );
  COND1XL U12242 ( .A(n17829), .B(n13434), .C(n11978), .Z(n13435) );
  CMX2X1 U12243 ( .A0(n13435), .A1(Poly2[28]), .S(n12211), .Z(n8982) );
  CIVX1 U12244 ( .A(Poly6[46]), .Z(n16956) );
  CEOX1 U12245 ( .A(Poly6[35]), .B(n16956), .Z(n13437) );
  CIVX2 U12246 ( .A(n13437), .Z(n13436) );
  CANR2X1 U12247 ( .A(n16063), .B(poly6_shifted[55]), .C(n13689), .D(n13436), 
        .Z(n13439) );
  COND4CX1 U12248 ( .A(n13437), .B(n13691), .C(n18219), .D(n13837), .Z(n13438)
         );
  CND2X1 U12249 ( .A(n13439), .B(n13438), .Z(n9648) );
  COND1XL U12250 ( .A(poly0_shifted[71]), .B(n18138), .C(n18137), .Z(n13441)
         );
  CMXI2X1 U12251 ( .A0(n13441), .A1(n13440), .S(n12291), .Z(n9506) );
  CIVX1 U12252 ( .A(poly6_shifted[17]), .Z(n13445) );
  CND3XL U12253 ( .A(n17718), .B(n13467), .C(n13452), .Z(n13442) );
  COND1XL U12254 ( .A(Poly6[53]), .B(n13467), .C(n13442), .Z(n13444) );
  CMXI2X1 U12255 ( .A0(n13445), .A1(n13444), .S(n16962), .Z(n9686) );
  CNR2XL U12256 ( .A(n17829), .B(Poly11[82]), .Z(n13504) );
  CIVDX2 U12257 ( .A(n13579), .Z0(n15843), .Z1(n13446) );
  COND4CX1 U12258 ( .A(Poly11[61]), .B(n13504), .C(n13028), .D(n13446), .Z(
        n13448) );
  CND2X1 U12259 ( .A(n15843), .B(Poly11[76]), .Z(n13447) );
  COND3X1 U12260 ( .A(Poly11[61]), .B(n13507), .C(n13448), .D(n13447), .Z(
        n11113) );
  COND1XL U12261 ( .A(Poly6[49]), .B(Poly6[38]), .C(n17705), .Z(n13451) );
  CMXI2X1 U12262 ( .A0(n12381), .A1(Poly6[48]), .S(n16063), .Z(n13450) );
  COND4CX1 U12263 ( .A(Poly6[38]), .B(Poly6[49]), .C(n13451), .D(n13450), .Z(
        n9645) );
  COND1XL U12264 ( .A(Poly12[115]), .B(Poly12[19]), .C(n17206), .Z(n13455) );
  CMXI2X1 U12265 ( .A0(n18053), .A1(Poly12[35]), .S(n12598), .Z(n13454) );
  COND4CX1 U12266 ( .A(Poly12[19]), .B(Poly12[115]), .C(n13455), .D(n13454), 
        .Z(n10497) );
  COND1XL U12267 ( .A(Poly12[122]), .B(Poly12[33]), .C(n18234), .Z(n13457) );
  CMXI2X1 U12268 ( .A0(n13522), .A1(poly12_shifted[65]), .S(n12598), .Z(n13456) );
  COND4CX1 U12269 ( .A(Poly12[33]), .B(Poly12[122]), .C(n13457), .D(n13456), 
        .Z(n10483) );
  CIVX2 U12270 ( .A(n15673), .Z(n16479) );
  COND1XL U12271 ( .A(Poly12[32]), .B(Poly12[121]), .C(n16479), .Z(n13459) );
  CMXI2X1 U12272 ( .A0(n18167), .A1(poly12_shifted[64]), .S(n12598), .Z(n13458) );
  COND4CX1 U12273 ( .A(Poly12[121]), .B(Poly12[32]), .C(n13459), .D(n13458), 
        .Z(n10484) );
  CND2X1 U12274 ( .A(n14292), .B(Poly12[17]), .Z(n13461) );
  CIVX1 U12275 ( .A(n17711), .Z(n14361) );
  CMXI2X1 U12276 ( .A0(n14361), .A1(Poly12[33]), .S(n12598), .Z(n13460) );
  COND3X1 U12277 ( .A(Poly12[17]), .B(n14295), .C(n13461), .D(n13460), .Z(
        n10499) );
  CMXI2X1 U12278 ( .A0(n13028), .A1(poly12_shifted[28]), .S(n12997), .Z(n13463) );
  CND2XL U12279 ( .A(n17755), .B(Poly12[123]), .Z(n13462) );
  CND2X1 U12280 ( .A(n13463), .B(n13462), .Z(n10520) );
  CIVX2 U12281 ( .A(n13467), .Z(n13681) );
  CANR2X1 U12282 ( .A(n16063), .B(Poly6[40]), .C(n13681), .D(Poly6[30]), .Z(
        n13466) );
  CIVXL U12283 ( .A(Poly6[30]), .Z(n13464) );
  COND4CX1 U12284 ( .A(n13683), .B(n13464), .C(n18142), .D(n13837), .Z(n13465)
         );
  CND2X1 U12285 ( .A(n13466), .B(n13465), .Z(n9653) );
  CND2X1 U12286 ( .A(n12068), .B(Poly2[69]), .Z(n16753) );
  CIVX1 U12287 ( .A(Poly2[69]), .Z(n13748) );
  CAN2X1 U12288 ( .A(n18234), .B(n13748), .Z(n13553) );
  COND1XL U12289 ( .A(Poly15[56]), .B(Poly15[30]), .C(n17063), .Z(n13470) );
  CMXI2X1 U12290 ( .A0(n18219), .A1(Poly15[45]), .S(n17376), .Z(n13469) );
  COND4CX1 U12291 ( .A(Poly15[30]), .B(Poly15[56]), .C(n13470), .D(n13469), 
        .Z(n9592) );
  CND2X1 U12292 ( .A(n17714), .B(Poly11[79]), .Z(n14190) );
  CIVXL U12293 ( .A(Poly11[79]), .Z(n13471) );
  CAN2X1 U12294 ( .A(n18017), .B(n13471), .Z(n13619) );
  CND2X1 U12295 ( .A(n13619), .B(Poly11[40]), .Z(n13473) );
  CMXI2X1 U12296 ( .A0(n11999), .A1(Poly11[55]), .S(n17683), .Z(n13472) );
  COND3X1 U12297 ( .A(Poly11[40]), .B(n14190), .C(n13473), .D(n13472), .Z(
        n11134) );
  CND2X1 U12298 ( .A(n15378), .B(poly5_shifted[67]), .Z(n13475) );
  CND2X1 U12299 ( .A(n17508), .B(poly5_shifted[53]), .Z(n13474) );
  COND3X1 U12300 ( .A(n15378), .B(n12006), .C(n13475), .D(n13474), .Z(n11473)
         );
  CEOXL U12301 ( .A(n16385), .B(dataselector[24]), .Z(n13476) );
  CENX1 U12302 ( .A(n17821), .B(n13476), .Z(n13477) );
  CANR1XL U12303 ( .A(n18234), .B(n13477), .C(n12003), .Z(n13478) );
  CMXI2X1 U12304 ( .A0(n13479), .A1(n13478), .S(n15799), .Z(n8764) );
  CND2X1 U12305 ( .A(n14310), .B(Poly6[4]), .Z(n13480) );
  COND4CX1 U12306 ( .A(n13481), .B(n12005), .C(n14310), .D(n13480), .Z(n9689)
         );
  CIVX2 U12307 ( .A(poly5_shifted[63]), .Z(n13502) );
  COND1XL U12308 ( .A(n17829), .B(n13502), .C(n13482), .Z(n13483) );
  CMX2X1 U12309 ( .A0(n13483), .A1(poly5_shifted[77]), .S(n15361), .Z(n11463)
         );
  CEOX1 U12310 ( .A(Poly6[37]), .B(n13833), .Z(n13485) );
  CIVX2 U12311 ( .A(n13485), .Z(n13484) );
  CANR2X1 U12312 ( .A(n16063), .B(Poly6[47]), .C(n13484), .D(n13681), .Z(
        n13487) );
  COND4CX1 U12313 ( .A(n13683), .B(n13485), .C(n18206), .D(n13837), .Z(n13486)
         );
  CND2X1 U12314 ( .A(n13487), .B(n13486), .Z(n9646) );
  CND2X1 U12315 ( .A(n17747), .B(Poly11[53]), .Z(n13490) );
  CMXI2X1 U12316 ( .A0(n16415), .A1(n13488), .S(Poly11[38]), .Z(n13489) );
  COND3X1 U12317 ( .A(n17683), .B(n12006), .C(n13490), .D(n13489), .Z(n11136)
         );
  CMXI2XL U12318 ( .A0(n16381), .A1(poly7_shifted[23]), .S(n17564), .Z(n13492)
         );
  CND2XL U12319 ( .A(n17545), .B(Poly7[410]), .Z(n13491) );
  CND2X1 U12320 ( .A(n13492), .B(n13491), .Z(n10093) );
  CND2X1 U12321 ( .A(n17755), .B(Poly6[52]), .Z(n13818) );
  COND4CXL U12322 ( .A(Poly6[41]), .B(n13815), .C(n18176), .D(n13837), .Z(
        n13495) );
  CND2XL U12323 ( .A(Poly6[51]), .B(n14166), .Z(n13494) );
  COND3X1 U12324 ( .A(Poly6[41]), .B(n13818), .C(n13495), .D(n13494), .Z(n9642) );
  CIVXL U12325 ( .A(Poly6[17]), .Z(n13497) );
  COND1XL U12326 ( .A(n13522), .B(poly6_shifted[17]), .C(n18193), .Z(n13496)
         );
  CMXI2X1 U12327 ( .A0(n13497), .A1(n13496), .S(n16962), .Z(n9676) );
  CMXI2XL U12328 ( .A0(n12013), .A1(Poly6[42]), .S(n14166), .Z(n13501) );
  CMXI2X1 U12329 ( .A0(n13499), .A1(n13498), .S(Poly6[32]), .Z(n13500) );
  CND2X1 U12330 ( .A(n13501), .B(n13500), .Z(n9651) );
  COND1XL U12331 ( .A(n13522), .B(poly5_shifted[49]), .C(n18193), .Z(n13503)
         );
  CMXI2X1 U12332 ( .A0(n13503), .A1(n13502), .S(n17935), .Z(n11477) );
  COND4CXL U12333 ( .A(Poly11[28]), .B(n13504), .C(n16381), .D(n11998), .Z(
        n13506) );
  CND2X1 U12334 ( .A(n17683), .B(Poly11[43]), .Z(n13505) );
  COND3X1 U12335 ( .A(Poly11[28]), .B(n13507), .C(n13506), .D(n13505), .Z(
        n11146) );
  COND1XL U12336 ( .A(Poly11[45]), .B(n13510), .C(n17714), .Z(n13509) );
  COND4CX1 U12337 ( .A(n13510), .B(Poly11[45]), .C(n13509), .D(n13508), .Z(
        n11129) );
  COND4CXL U12338 ( .A(Poly12[31]), .B(n14284), .C(n18206), .D(n13511), .Z(
        n13513) );
  CND2X1 U12339 ( .A(n12598), .B(poly12_shifted[63]), .Z(n13512) );
  COND3X1 U12340 ( .A(Poly12[31]), .B(n14287), .C(n13513), .D(n13512), .Z(
        n10485) );
  CND2X1 U12341 ( .A(n17930), .B(poly5_shifted[41]), .Z(n13515) );
  CND2X1 U12342 ( .A(n17545), .B(poly5_shifted[27]), .Z(n13514) );
  COND3X1 U12343 ( .A(n17932), .B(n17741), .C(n13515), .D(n13514), .Z(n11499)
         );
  CIVX2 U12344 ( .A(n15648), .Z(n17504) );
  CND2X1 U12345 ( .A(poly0_shifted[112]), .B(n17504), .Z(n13517) );
  COND2X1 U12346 ( .A(n16274), .B(Poly0[112]), .C(n15880), .D(n18167), .Z(
        n13516) );
  CND2X1 U12347 ( .A(n13517), .B(n13516), .Z(n9465) );
  CND2X1 U12348 ( .A(poly0_shifted[100]), .B(n16702), .Z(n13519) );
  COND2X1 U12349 ( .A(n16274), .B(poly0_shifted[118]), .C(n15880), .D(n12004), 
        .Z(n13518) );
  CND2X1 U12350 ( .A(n13519), .B(n13518), .Z(n9477) );
  CIVX2 U12351 ( .A(n15648), .Z(n17965) );
  CND2X1 U12352 ( .A(poly0_shifted[105]), .B(n17965), .Z(n13521) );
  COND2X1 U12353 ( .A(n16274), .B(Poly0[105]), .C(n15880), .D(n18189), .Z(
        n13520) );
  CND2X1 U12354 ( .A(n13521), .B(n13520), .Z(n9472) );
  CND2X1 U12355 ( .A(poly0_shifted[113]), .B(n17298), .Z(n13524) );
  COND2X1 U12356 ( .A(n16274), .B(Poly0[113]), .C(n15880), .D(n13522), .Z(
        n13523) );
  CND2X1 U12357 ( .A(n13524), .B(n13523), .Z(n9464) );
  CND2X1 U12358 ( .A(poly0_shifted[103]), .B(n17508), .Z(n13526) );
  COND2X1 U12359 ( .A(n16274), .B(Poly0[103]), .C(n15880), .D(n18138), .Z(
        n13525) );
  CND2X1 U12360 ( .A(n13526), .B(n13525), .Z(n9474) );
  CND2X1 U12361 ( .A(poly0_shifted[110]), .B(n17094), .Z(n13528) );
  COND2X1 U12362 ( .A(n16274), .B(Poly0[110]), .C(n15880), .D(n18160), .Z(
        n13527) );
  CND2X1 U12363 ( .A(n13528), .B(n13527), .Z(n9467) );
  CEOXL U12364 ( .A(Poly5[111]), .B(Poly5[124]), .Z(n13529) );
  CENX1 U12365 ( .A(Poly5[89]), .B(n13529), .Z(n13530) );
  COND2X1 U12366 ( .A(n13530), .B(n17744), .C(n13904), .D(n16939), .Z(n13531)
         );
  CAOR1X1 U12367 ( .A(poly5_shifted[117]), .B(n15403), .C(n13531), .Z(n11423)
         );
  CEOXL U12368 ( .A(Poly2[67]), .B(Poly2[27]), .Z(n13532) );
  CMXI2X1 U12369 ( .A0(n17364), .A1(n17366), .S(n13532), .Z(n13534) );
  CMXI2X1 U12370 ( .A0(n18138), .A1(Poly2[39]), .S(n12022), .Z(n13533) );
  CND2X1 U12371 ( .A(n13534), .B(n13533), .Z(n8971) );
  COND1XL U12372 ( .A(Poly1[342]), .B(Poly1[59]), .C(n18017), .Z(n13536) );
  CMXI2X1 U12373 ( .A0(n18116), .A1(poly1_shifted[81]), .S(n12012), .Z(n13535)
         );
  COND4CX1 U12374 ( .A(Poly1[59]), .B(Poly1[342]), .C(n13536), .D(n13535), .Z(
        n9287) );
  COND1XL U12375 ( .A(Poly1[338]), .B(Poly1[55]), .C(n17401), .Z(n13538) );
  CMXI2X1 U12376 ( .A0(n13428), .A1(poly1_shifted[77]), .S(n12012), .Z(n13537)
         );
  COND4CX1 U12377 ( .A(Poly1[55]), .B(Poly1[338]), .C(n13538), .D(n13537), .Z(
        n9291) );
  COND1XL U12378 ( .A(Poly1[346]), .B(Poly1[63]), .C(n17655), .Z(n13540) );
  CMXI2X1 U12379 ( .A0(n12013), .A1(poly1_shifted[85]), .S(n12012), .Z(n13539)
         );
  COND4CX1 U12380 ( .A(Poly1[63]), .B(Poly1[346]), .C(n13540), .D(n13539), .Z(
        n9283) );
  COND1XL U12381 ( .A(Poly1[337]), .B(Poly1[54]), .C(n17538), .Z(n13542) );
  CMXI2X1 U12382 ( .A0(n13812), .A1(poly1_shifted[76]), .S(n12012), .Z(n13541)
         );
  COND4CX1 U12383 ( .A(Poly1[54]), .B(Poly1[337]), .C(n13542), .D(n13541), .Z(
        n9292) );
  COND1XL U12384 ( .A(Poly1[53]), .B(Poly1[336]), .C(n17343), .Z(n13544) );
  CMXI2X1 U12385 ( .A0(n18108), .A1(poly1_shifted[75]), .S(n12012), .Z(n13543)
         );
  COND4CX1 U12386 ( .A(Poly1[336]), .B(Poly1[53]), .C(n13544), .D(n13543), .Z(
        n9293) );
  COND1XL U12387 ( .A(Poly5[86]), .B(Poly5[121]), .C(n17288), .Z(n13546) );
  CMXI2X1 U12388 ( .A0(n12004), .A1(Poly5[100]), .S(n12016), .Z(n13545) );
  COND4CX1 U12389 ( .A(Poly5[121]), .B(Poly5[86]), .C(n13546), .D(n13545), .Z(
        n11426) );
  COND1XL U12390 ( .A(Poly5[116]), .B(Poly5[94]), .C(n17705), .Z(n13548) );
  CMXI2X1 U12391 ( .A0(n13028), .A1(poly5_shifted[122]), .S(n12016), .Z(n13547) );
  COND4CX1 U12392 ( .A(Poly5[94]), .B(Poly5[116]), .C(n13548), .D(n13547), .Z(
        n11418) );
  COND1XL U12393 ( .A(Poly5[120]), .B(Poly5[98]), .C(n17634), .Z(n13550) );
  CMXI2X1 U12394 ( .A0(n18167), .A1(Poly5[112]), .S(n12016), .Z(n13549) );
  COND4CX1 U12395 ( .A(Poly5[98]), .B(Poly5[120]), .C(n13550), .D(n13549), .Z(
        n11414) );
  COND1XL U12396 ( .A(Poly6[4]), .B(Poly6[55]), .C(n18017), .Z(n13552) );
  CMXI2X1 U12397 ( .A0(n18160), .A1(Poly6[14]), .S(n13840), .Z(n13551) );
  COND4CX1 U12398 ( .A(Poly6[55]), .B(Poly6[4]), .C(n13552), .D(n13551), .Z(
        n9679) );
  CND2X1 U12399 ( .A(n12002), .B(n17826), .Z(n18188) );
  CND2X1 U12400 ( .A(n15361), .B(poly5_shifted[73]), .Z(n13555) );
  CND2X1 U12401 ( .A(n17755), .B(poly5_shifted[59]), .Z(n13554) );
  COND3X1 U12402 ( .A(n15361), .B(n17741), .C(n13555), .D(n13554), .Z(n11467)
         );
  CENX1 U12403 ( .A(dataselector[61]), .B(n18239), .Z(n13556) );
  CEOX1 U12404 ( .A(n13556), .B(dataselector[3]), .Z(n13557) );
  COND2XL U12405 ( .A(n13557), .B(n17495), .C(n12014), .D(n14944), .Z(n13558)
         );
  CAOR1X1 U12406 ( .A(n16410), .B(dataselector[10]), .C(n13558), .Z(n8785) );
  CND2X1 U12407 ( .A(n15361), .B(poly5_shifted[56]), .Z(n13560) );
  CND2X1 U12408 ( .A(n17705), .B(poly5_shifted[42]), .Z(n13559) );
  COND3X1 U12409 ( .A(n15361), .B(n12014), .C(n13560), .D(n13559), .Z(n11484)
         );
  COND1XL U12410 ( .A(Poly11[52]), .B(n13563), .C(n17714), .Z(n13562) );
  CMXI2X1 U12411 ( .A0(n18053), .A1(Poly11[67]), .S(n15843), .Z(n13561) );
  COND4CX1 U12412 ( .A(n13563), .B(Poly11[52]), .C(n13562), .D(n13561), .Z(
        n11122) );
  COND1XL U12413 ( .A(Poly13[519]), .B(Poly13[392]), .C(n17755), .Z(n13565) );
  CMXI2X1 U12414 ( .A0(n18034), .A1(poly13_shifted[420]), .S(n17043), .Z(
        n13564) );
  COND4CX1 U12415 ( .A(Poly13[392]), .B(Poly13[519]), .C(n13565), .D(n13564), 
        .Z(n10654) );
  COND1XL U12416 ( .A(Poly13[525]), .B(Poly13[398]), .C(n16700), .Z(n13567) );
  COND4CX1 U12417 ( .A(Poly13[398]), .B(Poly13[525]), .C(n13567), .D(n13566), 
        .Z(n10648) );
  COND1XL U12418 ( .A(Poly13[520]), .B(Poly13[393]), .C(n17094), .Z(n13569) );
  CMXI2X1 U12419 ( .A0(n11999), .A1(poly13_shifted[421]), .S(n17043), .Z(
        n13568) );
  COND4CX1 U12420 ( .A(Poly13[393]), .B(Poly13[520]), .C(n13569), .D(n13568), 
        .Z(n10653) );
  COND1XL U12421 ( .A(Poly13[514]), .B(Poly13[387]), .C(n17552), .Z(n13571) );
  CMXI2X1 U12422 ( .A0(n13522), .A1(poly13_shifted[415]), .S(n17043), .Z(
        n13570) );
  COND4CX1 U12423 ( .A(Poly13[387]), .B(Poly13[514]), .C(n13571), .D(n13570), 
        .Z(n10659) );
  CEOX1 U12424 ( .A(Poly10[31]), .B(Poly10[36]), .Z(n15951) );
  CMXI2XL U12425 ( .A0(n18228), .A1(poly10_shifted[41]), .S(n17962), .Z(n13575) );
  CENX1 U12426 ( .A(Poly10[38]), .B(Poly10[33]), .Z(n15905) );
  CENX1 U12427 ( .A(Poly10[17]), .B(n15905), .Z(n13573) );
  CND2X1 U12428 ( .A(n13573), .B(n16372), .Z(n13574) );
  CND2X1 U12429 ( .A(n13575), .B(n13574), .Z(n11074) );
  CMXI2XL U12430 ( .A0(n18105), .A1(poly10_shifted[42]), .S(n17962), .Z(n13578) );
  CENX1 U12431 ( .A(Poly10[39]), .B(Poly10[34]), .Z(n15941) );
  CENX1 U12432 ( .A(Poly10[18]), .B(n15941), .Z(n13576) );
  CND2X1 U12433 ( .A(n18047), .B(n13576), .Z(n13577) );
  CND2X1 U12434 ( .A(n13578), .B(n13577), .Z(n11073) );
  COND4CX1 U12435 ( .A(Poly11[49]), .B(n13619), .C(n12010), .D(n13446), .Z(
        n13581) );
  CND2X1 U12436 ( .A(n15843), .B(Poly11[64]), .Z(n13580) );
  COND3X1 U12437 ( .A(Poly11[49]), .B(n14190), .C(n13581), .D(n13580), .Z(
        n11125) );
  COND4CXL U12438 ( .A(Poly11[25]), .B(n13619), .C(n18142), .D(n11998), .Z(
        n13583) );
  CND2X1 U12439 ( .A(n17747), .B(Poly11[40]), .Z(n13582) );
  COND3X1 U12440 ( .A(Poly11[25]), .B(n14190), .C(n13583), .D(n13582), .Z(
        n11149) );
  COND1XL U12441 ( .A(Poly7[402]), .B(Poly7[22]), .C(n17535), .Z(n13585) );
  CMXI2X1 U12442 ( .A0(n13428), .A1(poly7_shifted[46]), .S(n12170), .Z(n13584)
         );
  COND4CX1 U12443 ( .A(Poly7[22]), .B(Poly7[402]), .C(n13585), .D(n13584), .Z(
        n10070) );
  CNR2X1 U12444 ( .A(n18116), .B(n17925), .Z(n13587) );
  CMXI2X1 U12445 ( .A0(n13587), .A1(Poly5[117]), .S(n13586), .Z(n13588) );
  CMX2X1 U12446 ( .A0(n13588), .A1(poly5_shifted[20]), .S(n17932), .Z(n11520)
         );
  CND2X1 U12447 ( .A(n15361), .B(poly5_shifted[75]), .Z(n13590) );
  CIVX2 U12448 ( .A(n15648), .Z(n17613) );
  CND2X1 U12449 ( .A(n17613), .B(poly5_shifted[61]), .Z(n13589) );
  COND3X1 U12450 ( .A(n17935), .B(n17185), .C(n13590), .D(n13589), .Z(n11465)
         );
  CIVXL U12451 ( .A(Poly5[114]), .Z(n13591) );
  CIVXL U12452 ( .A(Poly1[344]), .Z(n13592) );
  CIVXL U12453 ( .A(Poly6[44]), .Z(n13593) );
  CND2X1 U12454 ( .A(n13593), .B(n13833), .Z(n13594) );
  CND2X1 U12455 ( .A(n16323), .B(n13594), .Z(n13596) );
  CMXI2X1 U12456 ( .A0(n18034), .A1(Poly6[54]), .S(n16063), .Z(n13595) );
  COND4CX1 U12457 ( .A(Poly6[44]), .B(Poly6[55]), .C(n13596), .D(n13595), .Z(
        n9639) );
  CEOXL U12458 ( .A(Poly12[28]), .B(Poly12[117]), .Z(n13599) );
  COND1XL U12459 ( .A(Poly12[124]), .B(n13599), .C(n16702), .Z(n13598) );
  CMXI2X1 U12460 ( .A0(n13028), .A1(poly12_shifted[60]), .S(n12598), .Z(n13597) );
  COND4CX1 U12461 ( .A(n13599), .B(Poly12[124]), .C(n13598), .D(n13597), .Z(
        n10488) );
  CIVX2 U12462 ( .A(n15648), .Z(n17285) );
  COND1XL U12463 ( .A(Poly12[16]), .B(Poly12[112]), .C(n17285), .Z(n13601) );
  CMXI2X1 U12464 ( .A0(n12010), .A1(Poly12[32]), .S(n12598), .Z(n13600) );
  COND4CX1 U12465 ( .A(Poly12[112]), .B(Poly12[16]), .C(n13601), .D(n13600), 
        .Z(n10500) );
  CEOX1 U12466 ( .A(Poly12[27]), .B(Poly12[123]), .Z(n13602) );
  CEOXL U12467 ( .A(Poly12[120]), .B(Poly12[24]), .Z(n13605) );
  CND2X1 U12468 ( .A(n14292), .B(n13605), .Z(n13604) );
  CMXI2X1 U12469 ( .A0(n18142), .A1(poly12_shifted[56]), .S(n12598), .Z(n13603) );
  COND3X1 U12470 ( .A(n13605), .B(n14295), .C(n13604), .D(n13603), .Z(n10492)
         );
  COND1XL U12471 ( .A(Poly13[521]), .B(Poly13[162]), .C(n17401), .Z(n13607) );
  CMXI2X1 U12472 ( .A0(n18167), .A1(poly13_shifted[190]), .S(n13014), .Z(
        n13606) );
  COND4CX1 U12473 ( .A(Poly13[162]), .B(Poly13[521]), .C(n13607), .D(n13606), 
        .Z(n10884) );
  COND1XL U12474 ( .A(Poly13[522]), .B(Poly13[163]), .C(n17362), .Z(n13609) );
  CMXI2X1 U12475 ( .A0(n13522), .A1(poly13_shifted[191]), .S(n13014), .Z(
        n13608) );
  COND4CX1 U12476 ( .A(Poly13[163]), .B(Poly13[522]), .C(n13609), .D(n13608), 
        .Z(n10883) );
  COND1XL U12477 ( .A(Poly11[51]), .B(n13612), .C(n17714), .Z(n13611) );
  CMXI2X1 U12478 ( .A0(n13428), .A1(Poly11[66]), .S(n15843), .Z(n13610) );
  COND4CX1 U12479 ( .A(n13612), .B(Poly11[51]), .C(n13611), .D(n13610), .Z(
        n11123) );
  COND1XL U12480 ( .A(Poly0[210]), .B(Poly0[158]), .C(n17705), .Z(n13614) );
  CANR2X1 U12481 ( .A(n18167), .B(n15960), .C(poly0_shifted[194]), .D(n17314), 
        .Z(n13613) );
  COND4CX1 U12482 ( .A(Poly0[158]), .B(Poly0[210]), .C(n13614), .D(n13613), 
        .Z(n9401) );
  COND1XL U12483 ( .A(Poly0[218]), .B(Poly0[166]), .C(n17466), .Z(n13616) );
  CANR2X1 U12484 ( .A(n13994), .B(n15960), .C(poly0_shifted[202]), .D(n15671), 
        .Z(n13615) );
  COND4CX1 U12485 ( .A(Poly0[166]), .B(Poly0[218]), .C(n13616), .D(n13615), 
        .Z(n9393) );
  COND1XL U12486 ( .A(Poly0[216]), .B(Poly0[164]), .C(n18017), .Z(n13618) );
  CANR2X1 U12487 ( .A(n18034), .B(n15960), .C(poly0_shifted[200]), .D(n15671), 
        .Z(n13617) );
  COND4CX1 U12488 ( .A(Poly0[164]), .B(Poly0[216]), .C(n13618), .D(n13617), 
        .Z(n9395) );
  CND2X1 U12489 ( .A(n13619), .B(Poly11[58]), .Z(n13621) );
  CMXI2X1 U12490 ( .A0(n18189), .A1(Poly11[73]), .S(n15843), .Z(n13620) );
  COND3X1 U12491 ( .A(Poly11[58]), .B(n14190), .C(n13621), .D(n13620), .Z(
        n11116) );
  COND1XL U12492 ( .A(Poly0[215]), .B(Poly0[163]), .C(n18234), .Z(n13623) );
  CANR2X1 U12493 ( .A(n18241), .B(n15960), .C(poly0_shifted[199]), .D(n17314), 
        .Z(n13622) );
  COND4CX1 U12494 ( .A(Poly0[163]), .B(Poly0[215]), .C(n13623), .D(n13622), 
        .Z(n9396) );
  COND1XL U12495 ( .A(Poly0[211]), .B(Poly0[159]), .C(n17755), .Z(n13625) );
  CANR2X1 U12496 ( .A(n14297), .B(n15960), .C(poly0_shifted[195]), .D(n17314), 
        .Z(n13624) );
  COND4CX1 U12497 ( .A(Poly0[159]), .B(Poly0[211]), .C(n13625), .D(n13624), 
        .Z(n9400) );
  CIVX2 U12498 ( .A(n15673), .Z(n17121) );
  COND1XL U12499 ( .A(Poly6[49]), .B(Poly6[31]), .C(n17121), .Z(n13627) );
  CMXI2X1 U12500 ( .A0(n18189), .A1(Poly6[41]), .S(n14166), .Z(n13626) );
  COND4CX1 U12501 ( .A(Poly6[31]), .B(Poly6[49]), .C(n13627), .D(n13626), .Z(
        n9652) );
  COND1XL U12502 ( .A(Poly6[28]), .B(Poly6[46]), .C(n16312), .Z(n13629) );
  CMXI2X1 U12503 ( .A0(n14754), .A1(Poly6[38]), .S(n14166), .Z(n13628) );
  COND4CX1 U12504 ( .A(Poly6[46]), .B(Poly6[28]), .C(n13629), .D(n13628), .Z(
        n9655) );
  CND2X1 U12505 ( .A(n13815), .B(Poly6[24]), .Z(n13631) );
  CMXI2X1 U12506 ( .A0(n13428), .A1(Poly6[34]), .S(n14166), .Z(n13630) );
  COND3X1 U12507 ( .A(Poly6[24]), .B(n13818), .C(n13631), .D(n13630), .Z(n9659) );
  CND2X1 U12508 ( .A(n13815), .B(Poly6[34]), .Z(n13633) );
  CMXI2X1 U12509 ( .A0(n13028), .A1(Poly6[44]), .S(n14166), .Z(n13632) );
  COND3X1 U12510 ( .A(Poly6[34]), .B(n13818), .C(n13633), .D(n13632), .Z(n9649) );
  CND2X1 U12511 ( .A(n16961), .B(Poly6[26]), .Z(n13635) );
  CMXI2X1 U12512 ( .A0(n12004), .A1(Poly6[36]), .S(n14166), .Z(n13634) );
  COND3X1 U12513 ( .A(Poly6[26]), .B(n16957), .C(n13635), .D(n13634), .Z(n9657) );
  CEOX1 U12514 ( .A(n18239), .B(dataselector[62]), .Z(n16135) );
  CEOX1 U12515 ( .A(dataselector[11]), .B(n16135), .Z(n13636) );
  CANR2X1 U12516 ( .A(n16410), .B(dataselector[18]), .C(n17523), .D(n13636), 
        .Z(n13638) );
  CND2XL U12517 ( .A(n18210), .B(n17832), .Z(n13637) );
  CND2X1 U12518 ( .A(n13638), .B(n13637), .Z(n8777) );
  CENX1 U12519 ( .A(dataselector[58]), .B(n18239), .Z(n15645) );
  CENX1 U12520 ( .A(n14017), .B(n15645), .Z(n15919) );
  COND1XL U12521 ( .A(dataselector[9]), .B(n15919), .C(n17535), .Z(n13640) );
  CANR2X1 U12522 ( .A(n12381), .B(n17832), .C(dataselector[16]), .D(n16410), 
        .Z(n13639) );
  COND4CX1 U12523 ( .A(n15919), .B(dataselector[9]), .C(n13640), .D(n13639), 
        .Z(n8779) );
  CEOXL U12524 ( .A(Poly0[204]), .B(Poly0[152]), .Z(n13641) );
  CND2XL U12525 ( .A(n17356), .B(n13641), .Z(n13643) );
  CND2X1 U12526 ( .A(n17314), .B(poly0_shifted[188]), .Z(n13642) );
  COND4CX1 U12527 ( .A(n12014), .B(n13643), .C(n15671), .D(n13642), .Z(n9407)
         );
  CIVXL U12528 ( .A(n17711), .Z(n14716) );
  CMXI2X1 U12529 ( .A0(n14716), .A1(Poly6[1]), .S(n14310), .Z(n13644) );
  CIVX2 U12530 ( .A(n15648), .Z(n17280) );
  CND2X1 U12531 ( .A(n17280), .B(Poly6[47]), .Z(n13864) );
  CND2X1 U12532 ( .A(n13644), .B(n13864), .Z(n9692) );
  CMXI2X1 U12533 ( .A0(n17313), .A1(n13647), .S(Poly2[34]), .Z(n13646) );
  CMXI2X1 U12534 ( .A0(n18160), .A1(Poly2[46]), .S(n17306), .Z(n13645) );
  CND2X1 U12535 ( .A(n13646), .B(n13645), .Z(n8964) );
  CMXI2X1 U12536 ( .A0(n17313), .A1(n13647), .S(Poly2[21]), .Z(n13649) );
  CMXI2X1 U12537 ( .A0(n14361), .A1(Poly2[33]), .S(n17306), .Z(n13648) );
  CND2X1 U12538 ( .A(n13649), .B(n13648), .Z(n8977) );
  CND2X1 U12539 ( .A(n13815), .B(Poly6[1]), .Z(n13651) );
  CMXI2X1 U12540 ( .A0(n16381), .A1(Poly6[11]), .S(n14310), .Z(n13650) );
  COND3X1 U12541 ( .A(Poly6[1]), .B(n13818), .C(n13651), .D(n13650), .Z(n9682)
         );
  COND1XL U12542 ( .A(Poly0[205]), .B(Poly0[153]), .C(n17755), .Z(n13653) );
  CANR2X1 U12543 ( .A(n16381), .B(n15960), .C(n15671), .D(poly0_shifted[189]), 
        .Z(n13652) );
  COND4CX1 U12544 ( .A(Poly0[153]), .B(Poly0[205]), .C(n13653), .D(n13652), 
        .Z(n9406) );
  COND1XL U12545 ( .A(Poly0[203]), .B(Poly0[151]), .C(n17533), .Z(n13655) );
  CANR2X1 U12546 ( .A(n18189), .B(n15960), .C(n15671), .D(poly0_shifted[187]), 
        .Z(n13654) );
  COND4CX1 U12547 ( .A(Poly0[151]), .B(Poly0[203]), .C(n13655), .D(n13654), 
        .Z(n9408) );
  COND1XL U12548 ( .A(Poly0[206]), .B(Poly0[154]), .C(n17634), .Z(n13657) );
  CANR2X1 U12549 ( .A(n13028), .B(n15960), .C(n17314), .D(poly0_shifted[190]), 
        .Z(n13656) );
  COND4CX1 U12550 ( .A(Poly0[154]), .B(Poly0[206]), .C(n13657), .D(n13656), 
        .Z(n9405) );
  COND1XL U12551 ( .A(Poly0[207]), .B(Poly0[155]), .C(n16919), .Z(n13659) );
  CANR2X1 U12552 ( .A(n18219), .B(n15960), .C(n17314), .D(poly0_shifted[191]), 
        .Z(n13658) );
  COND4CX1 U12553 ( .A(Poly0[155]), .B(Poly0[207]), .C(n13659), .D(n13658), 
        .Z(n9404) );
  CND2X1 U12554 ( .A(n16695), .B(Poly8[82]), .Z(n13875) );
  CIVXL U12555 ( .A(Poly8[67]), .Z(n13661) );
  CANR4CXL U12556 ( .A(Poly8[82]), .B(n13661), .C(n17076), .D(n13660), .Z(
        n13662) );
  CND2XL U12557 ( .A(n13663), .B(n13662), .Z(n13665) );
  CND2X1 U12558 ( .A(n17750), .B(poly8_shifted[95]), .Z(n13664) );
  COND3X1 U12559 ( .A(Poly8[67]), .B(n13875), .C(n13665), .D(n13664), .Z(
        n11320) );
  CIVXL U12560 ( .A(Poly8[82]), .Z(n13666) );
  CND2IXL U12561 ( .B(n17160), .A(n13666), .Z(n13667) );
  CIVX2 U12562 ( .A(n13667), .Z(n13872) );
  CIVXL U12563 ( .A(n12175), .Z(n13668) );
  COND4CX1 U12564 ( .A(Poly8[1]), .B(n13872), .C(n18206), .D(n13668), .Z(
        n13670) );
  CND2X1 U12565 ( .A(n12175), .B(Poly8[15]), .Z(n13669) );
  COND3X1 U12566 ( .A(Poly8[1]), .B(n13875), .C(n13670), .D(n13669), .Z(n11386) );
  COND1XL U12567 ( .A(Poly5[97]), .B(Poly5[119]), .C(n17362), .Z(n13672) );
  CMXI2X1 U12568 ( .A0(n18206), .A1(Poly5[111]), .S(n12016), .Z(n13671) );
  COND4CX1 U12569 ( .A(Poly5[119]), .B(Poly5[97]), .C(n13672), .D(n13671), .Z(
        n11415) );
  COND1XL U12570 ( .A(Poly5[122]), .B(Poly5[87]), .C(n17280), .Z(n13674) );
  CMXI2X1 U12571 ( .A0(n11994), .A1(Poly5[101]), .S(n15403), .Z(n13673) );
  COND4CX1 U12572 ( .A(Poly5[87]), .B(Poly5[122]), .C(n13674), .D(n13673), .Z(
        n11425) );
  CMXI2X1 U12573 ( .A0(n16381), .A1(poly12_shifted[27]), .S(n12997), .Z(n13676) );
  CND2X1 U12574 ( .A(n17613), .B(Poly12[122]), .Z(n13675) );
  CND2X1 U12575 ( .A(n13676), .B(n13675), .Z(n10521) );
  CMXI2X1 U12576 ( .A0(n16381), .A1(poly3_shifted[25]), .S(n15737), .Z(n13678)
         );
  CND2X1 U12577 ( .A(n17343), .B(Poly3[81]), .Z(n13677) );
  CND2X1 U12578 ( .A(n13678), .B(n13677), .Z(n8929) );
  COND1XL U12579 ( .A(poly0_shifted[69]), .B(n11990), .C(n18134), .Z(n13680)
         );
  CMXI2X1 U12580 ( .A0(n13680), .A1(n13679), .S(n12291), .Z(n9508) );
  CANR2X1 U12581 ( .A(n14310), .B(Poly6[30]), .C(n13681), .D(Poly6[20]), .Z(
        n13685) );
  CIVXL U12582 ( .A(Poly6[20]), .Z(n13682) );
  COND4CXL U12583 ( .A(n13683), .B(n13682), .C(n18105), .D(n16962), .Z(n13684)
         );
  CND2X1 U12584 ( .A(n13685), .B(n13684), .Z(n9663) );
  CANR2X1 U12585 ( .A(n13840), .B(Poly6[12]), .C(Poly6[2]), .D(n13689), .Z(
        n13688) );
  COND4CX1 U12586 ( .A(n13691), .B(n13686), .C(n13028), .D(n16962), .Z(n13687)
         );
  CND2X1 U12587 ( .A(n13688), .B(n13687), .Z(n9681) );
  CANR2X1 U12588 ( .A(n16063), .B(Poly6[52]), .C(n13689), .D(Poly6[42]), .Z(
        n13693) );
  CIVXL U12589 ( .A(Poly6[42]), .Z(n13690) );
  COND4CX1 U12590 ( .A(n13691), .B(n13690), .C(n18082), .D(n13837), .Z(n13692)
         );
  CND2X1 U12591 ( .A(n13693), .B(n13692), .Z(n9641) );
  COND1XL U12592 ( .A(Poly0[103]), .B(Poly0[202]), .C(n17714), .Z(n13695) );
  CANR2X1 U12593 ( .A(n15880), .B(poly0_shifted[139]), .C(n18249), .D(n16274), 
        .Z(n13694) );
  COND4CX1 U12594 ( .A(Poly0[202]), .B(Poly0[103]), .C(n13695), .D(n13694), 
        .Z(n9456) );
  COND1XL U12595 ( .A(Poly0[205]), .B(Poly0[106]), .C(n17714), .Z(n13697) );
  COND4CX1 U12596 ( .A(Poly0[106]), .B(Poly0[205]), .C(n13697), .D(n13696), 
        .Z(n9453) );
  COND1XL U12597 ( .A(Poly5[121]), .B(Poly5[1]), .C(n17245), .Z(n13699) );
  CMXI2X1 U12598 ( .A0(n18206), .A1(poly5_shifted[29]), .S(n17932), .Z(n13698)
         );
  COND4CX1 U12599 ( .A(Poly5[1]), .B(Poly5[121]), .C(n13699), .D(n13698), .Z(
        n11511) );
  COND1XL U12600 ( .A(Poly5[119]), .B(Poly5[124]), .C(n16644), .Z(n13701) );
  CMXI2X1 U12601 ( .A0(n18219), .A1(poly5_shifted[27]), .S(n17932), .Z(n13700)
         );
  COND4CX1 U12602 ( .A(Poly5[124]), .B(Poly5[119]), .C(n13701), .D(n13700), 
        .Z(n11513) );
  CIVX2 U12603 ( .A(n17259), .Z(n17158) );
  COND1XL U12604 ( .A(Poly2[37]), .B(Poly2[64]), .C(n17158), .Z(n13703) );
  CIVXL U12605 ( .A(n17076), .Z(n14297) );
  CMXI2X1 U12606 ( .A0(n14297), .A1(Poly2[49]), .S(n17306), .Z(n13702) );
  COND4CX1 U12607 ( .A(Poly2[64]), .B(Poly2[37]), .C(n13703), .D(n13702), .Z(
        n8961) );
  CEOXL U12608 ( .A(Poly3[73]), .B(Poly3[48]), .Z(n13706) );
  COND1XL U12609 ( .A(Poly3[81]), .B(n13706), .C(n16479), .Z(n13705) );
  CMXI2X1 U12610 ( .A0(n18105), .A1(poly3_shifted[76]), .S(n17262), .Z(n13704)
         );
  COND4CX1 U12611 ( .A(n13706), .B(Poly3[81]), .C(n13705), .D(n13704), .Z(
        n8878) );
  CIVX2 U12612 ( .A(n17259), .Z(n17390) );
  COND1XL U12613 ( .A(Poly5[122]), .B(Poly5[2]), .C(n17390), .Z(n13708) );
  CMXI2X1 U12614 ( .A0(n18167), .A1(poly5_shifted[30]), .S(n17930), .Z(n13707)
         );
  COND4CX1 U12615 ( .A(Poly5[2]), .B(Poly5[122]), .C(n13708), .D(n13707), .Z(
        n11510) );
  COND1XL U12616 ( .A(Poly5[3]), .B(Poly5[123]), .C(n17598), .Z(n13710) );
  CMXI2X1 U12617 ( .A0(n18048), .A1(poly5_shifted[31]), .S(n17932), .Z(n13709)
         );
  COND4CX1 U12618 ( .A(Poly5[123]), .B(Poly5[3]), .C(n13710), .D(n13709), .Z(
        n11509) );
  COND1XL U12619 ( .A(Poly5[0]), .B(Poly5[120]), .C(n17295), .Z(n13712) );
  CMXI2X1 U12620 ( .A0(n18160), .A1(poly5_shifted[28]), .S(n17930), .Z(n13711)
         );
  COND4CX1 U12621 ( .A(Poly5[120]), .B(Poly5[0]), .C(n13712), .D(n13711), .Z(
        n11512) );
  CIVX2 U12622 ( .A(n15673), .Z(n17198) );
  COND1XL U12623 ( .A(Poly1[337]), .B(Poly1[21]), .C(n17198), .Z(n13714) );
  CMXI2X1 U12624 ( .A0(n12010), .A1(poly1_shifted[43]), .S(n12299), .Z(n13713)
         );
  COND4CX1 U12625 ( .A(Poly1[21]), .B(Poly1[337]), .C(n13714), .D(n13713), .Z(
        n9325) );
  COND1XL U12626 ( .A(Poly1[338]), .B(Poly1[22]), .C(n18234), .Z(n13716) );
  CMXI2X1 U12627 ( .A0(n14765), .A1(poly1_shifted[44]), .S(n12299), .Z(n13715)
         );
  COND4CX1 U12628 ( .A(Poly1[22]), .B(Poly1[338]), .C(n13716), .D(n13715), .Z(
        n9324) );
  CIVX1 U12629 ( .A(Poly1[341]), .Z(n14356) );
  CND2X1 U12630 ( .A(n14356), .B(n13717), .Z(n13718) );
  CND2X1 U12631 ( .A(n16323), .B(n13718), .Z(n13720) );
  CMXI2X1 U12632 ( .A0(n12004), .A1(poly1_shifted[47]), .S(n12299), .Z(n13719)
         );
  COND4CX1 U12633 ( .A(Poly1[25]), .B(Poly1[341]), .C(n13720), .D(n13719), .Z(
        n9321) );
  COND1XL U12634 ( .A(Poly1[345]), .B(Poly1[29]), .C(n17705), .Z(n13722) );
  CMXI2X1 U12635 ( .A0(n18142), .A1(poly1_shifted[51]), .S(n12299), .Z(n13721)
         );
  COND4CX1 U12636 ( .A(Poly1[29]), .B(Poly1[345]), .C(n13722), .D(n13721), .Z(
        n9317) );
  COND1XL U12637 ( .A(Poly1[343]), .B(Poly1[27]), .C(n17755), .Z(n13724) );
  CMXI2X1 U12638 ( .A0(n14754), .A1(poly1_shifted[49]), .S(n12299), .Z(n13723)
         );
  COND4CX1 U12639 ( .A(Poly1[27]), .B(Poly1[343]), .C(n13724), .D(n13723), .Z(
        n9319) );
  COND1XL U12640 ( .A(Poly1[344]), .B(Poly1[28]), .C(n17072), .Z(n13726) );
  CMXI2X1 U12641 ( .A0(n18138), .A1(poly1_shifted[50]), .S(n12299), .Z(n13725)
         );
  COND4CX1 U12642 ( .A(Poly1[28]), .B(Poly1[344]), .C(n13726), .D(n13725), .Z(
        n9318) );
  COND1XL U12643 ( .A(Poly1[342]), .B(Poly1[26]), .C(n18017), .Z(n13728) );
  CMXI2X1 U12644 ( .A0(n11984), .A1(poly1_shifted[48]), .S(n12299), .Z(n13727)
         );
  COND4CX1 U12645 ( .A(Poly1[26]), .B(Poly1[342]), .C(n13728), .D(n13727), .Z(
        n9320) );
  CANR2X1 U12646 ( .A(n12010), .B(n17832), .C(dataselector[0]), .D(n16410), 
        .Z(n13730) );
  CND2X1 U12647 ( .A(n13730), .B(n13729), .Z(n8795) );
  CENX1 U12648 ( .A(Poly10[37]), .B(n13731), .Z(n15942) );
  COND1XL U12649 ( .A(Poly10[16]), .B(n15942), .C(n17136), .Z(n13733) );
  COND4CX1 U12650 ( .A(n15942), .B(Poly10[16]), .C(n13733), .D(n13732), .Z(
        n11075) );
  COND1XL U12651 ( .A(Poly10[34]), .B(Poly10[13]), .C(n16427), .Z(n13735) );
  CMXI2X1 U12652 ( .A0(n18249), .A1(Poly10[25]), .S(n17962), .Z(n13734) );
  COND4CX1 U12653 ( .A(Poly10[13]), .B(Poly10[34]), .C(n13735), .D(n13734), 
        .Z(n11078) );
  COND1XL U12654 ( .A(Poly10[4]), .B(Poly10[42]), .C(n17178), .Z(n13737) );
  CMXI2X1 U12655 ( .A0(n18167), .A1(Poly10[16]), .S(n17962), .Z(n13736) );
  COND4CX1 U12656 ( .A(Poly10[42]), .B(Poly10[4]), .C(n13737), .D(n13736), .Z(
        n11087) );
  COND1XL U12657 ( .A(Poly10[10]), .B(Poly10[31]), .C(n17538), .Z(n13739) );
  CMXI2X1 U12658 ( .A0(n14487), .A1(Poly10[22]), .S(n17962), .Z(n13738) );
  COND4CX1 U12659 ( .A(Poly10[31]), .B(Poly10[10]), .C(n13739), .D(n13738), 
        .Z(n11081) );
  COND1XL U12660 ( .A(Poly12[123]), .B(Poly12[34]), .C(n18234), .Z(n13741) );
  CMXI2X1 U12661 ( .A0(n18210), .A1(poly12_shifted[66]), .S(n12598), .Z(n13740) );
  COND4CX1 U12662 ( .A(Poly12[34]), .B(Poly12[123]), .C(n13741), .D(n13740), 
        .Z(n10482) );
  COND1XL U12663 ( .A(Poly5[4]), .B(Poly5[124]), .C(n17527), .Z(n13743) );
  CMXI2X1 U12664 ( .A0(n18210), .A1(poly5_shifted[32]), .S(n17932), .Z(n13742)
         );
  COND4CX1 U12665 ( .A(Poly5[124]), .B(Poly5[4]), .C(n13743), .D(n13742), .Z(
        n11508) );
  COND1XL U12666 ( .A(Poly5[122]), .B(Poly5[100]), .C(n17401), .Z(n13745) );
  CMXI2X1 U12667 ( .A0(n18210), .A1(Poly5[114]), .S(n13904), .Z(n13744) );
  COND4CX1 U12668 ( .A(Poly5[100]), .B(Poly5[122]), .C(n13745), .D(n13744), 
        .Z(n11412) );
  COND1XL U12669 ( .A(Poly13[523]), .B(Poly13[164]), .C(n17634), .Z(n13747) );
  CMXI2X1 U12670 ( .A0(n18210), .A1(poly13_shifted[192]), .S(n13014), .Z(
        n13746) );
  COND4CX1 U12671 ( .A(Poly13[164]), .B(Poly13[523]), .C(n13747), .D(n13746), 
        .Z(n10882) );
  CND2X1 U12672 ( .A(Poly2[29]), .B(n13748), .Z(n13755) );
  CNR2X1 U12673 ( .A(Poly2[29]), .B(n13748), .Z(n13751) );
  CIVX2 U12674 ( .A(n13754), .Z(n14773) );
  CIVX1 U12675 ( .A(n14772), .Z(n16750) );
  CND2X1 U12676 ( .A(n13755), .B(n16750), .Z(n13749) );
  COND1XL U12677 ( .A(n13751), .B(n13749), .C(n12002), .Z(n13750) );
  COND4CX1 U12678 ( .A(n13751), .B(n14773), .C(n13750), .D(n12021), .Z(n13753)
         );
  CND2X1 U12679 ( .A(n12022), .B(Poly2[41]), .Z(n13752) );
  COND3X1 U12680 ( .A(n13755), .B(n13754), .C(n13753), .D(n13752), .Z(n8969)
         );
  COND1XL U12681 ( .A(Poly10[12]), .B(n13756), .C(n17721), .Z(n13757) );
  CMXI2X1 U12682 ( .A0(n13757), .A1(Poly10[24]), .S(n17962), .Z(n13758) );
  COND11X1 U12683 ( .A(Poly10[33]), .B(n17829), .C(n13759), .D(n13758), .Z(
        n11079) );
  CMXI2X1 U12684 ( .A0(n18138), .A1(poly12_shifted[23]), .S(n12997), .Z(n13760) );
  CND2X1 U12685 ( .A(n13760), .B(n14110), .Z(n10525) );
  COND1XL U12686 ( .A(Poly6[49]), .B(Poly6[13]), .C(n16326), .Z(n13762) );
  CMXI2X1 U12687 ( .A0(n11999), .A1(Poly6[23]), .S(n14310), .Z(n13761) );
  COND4CX1 U12688 ( .A(Poly6[13]), .B(Poly6[49]), .C(n13762), .D(n13761), .Z(
        n9670) );
  COND1XL U12689 ( .A(Poly9[107]), .B(Poly9[86]), .C(n17298), .Z(n13764) );
  CIVXL U12690 ( .A(n17711), .Z(n13812) );
  CMXI2X1 U12691 ( .A0(n13812), .A1(poly9_shifted[108]), .S(n12262), .Z(n13763) );
  COND4CX1 U12692 ( .A(Poly9[86]), .B(Poly9[107]), .C(n13764), .D(n13763), .Z(
        n11208) );
  CND2X1 U12693 ( .A(n15737), .B(poly3_shifted[15]), .Z(n13765) );
  COND4CX1 U12694 ( .A(n16950), .B(n13766), .C(n15737), .D(n13765), .Z(n8939)
         );
  CND2X1 U12695 ( .A(n12185), .B(poly11_shifted[22]), .Z(n13767) );
  COND3X1 U12696 ( .A(n12185), .B(n17718), .C(n13767), .D(n14303), .Z(n11182)
         );
  CIVX2 U12697 ( .A(n15648), .Z(n17998) );
  COND1XL U12698 ( .A(Poly1[342]), .B(Poly1[204]), .C(n17998), .Z(n13769) );
  CMXI2X1 U12699 ( .A0(n11999), .A1(poly1_shifted[226]), .S(n17053), .Z(n13768) );
  COND4CX1 U12700 ( .A(Poly1[204]), .B(Poly1[342]), .C(n13769), .D(n13768), 
        .Z(n9142) );
  COND1XL U12701 ( .A(Poly1[340]), .B(Poly1[57]), .C(n18047), .Z(n13771) );
  CMXI2X1 U12702 ( .A0(n12004), .A1(poly1_shifted[79]), .S(n12012), .Z(n13770)
         );
  COND4CX1 U12703 ( .A(Poly1[57]), .B(Poly1[340]), .C(n13771), .D(n13770), .Z(
        n9289) );
  COND1XL U12704 ( .A(Poly5[118]), .B(Poly5[96]), .C(n17144), .Z(n13773) );
  CMXI2X1 U12705 ( .A0(n18160), .A1(poly5_shifted[124]), .S(n13904), .Z(n13772) );
  COND4CX1 U12706 ( .A(Poly5[96]), .B(Poly5[118]), .C(n13773), .D(n13772), .Z(
        n11416) );
  COND1XL U12707 ( .A(Poly5[121]), .B(Poly5[99]), .C(n17488), .Z(n13775) );
  CMXI2X1 U12708 ( .A0(n18048), .A1(Poly5[113]), .S(n12016), .Z(n13774) );
  COND4CX1 U12709 ( .A(Poly5[99]), .B(Poly5[121]), .C(n13775), .D(n13774), .Z(
        n11413) );
  COND1XL U12710 ( .A(Poly1[344]), .B(Poly1[206]), .C(n17356), .Z(n13777) );
  CMXI2X1 U12711 ( .A0(n18249), .A1(poly1_shifted[228]), .S(n17053), .Z(n13776) );
  COND4CX1 U12712 ( .A(Poly1[206]), .B(Poly1[344]), .C(n13777), .D(n13776), 
        .Z(n9140) );
  COND1XL U12713 ( .A(Poly1[336]), .B(Poly1[198]), .C(n16695), .Z(n13779) );
  CMXI2X1 U12714 ( .A0(n18048), .A1(poly1_shifted[220]), .S(n17053), .Z(n13778) );
  COND4CX1 U12715 ( .A(Poly1[198]), .B(Poly1[336]), .C(n13779), .D(n13778), 
        .Z(n9148) );
  CEOX1 U12716 ( .A(n14017), .B(dataselector[59]), .Z(n14448) );
  COND1XL U12717 ( .A(n11999), .B(n13783), .C(n13782), .Z(n13785) );
  CND2X1 U12718 ( .A(n17634), .B(Poly10[11]), .Z(n13784) );
  CMXI2X1 U12719 ( .A0(Poly10[32]), .A1(n13785), .S(n13784), .Z(n13786) );
  CAOR1X1 U12720 ( .A(Poly10[23]), .B(n17962), .C(n13786), .Z(n11080) );
  CND2X1 U12721 ( .A(n17731), .B(poly9_shifted[18]), .Z(n13788) );
  CND2X1 U12722 ( .A(n17072), .B(Poly9[112]), .Z(n13787) );
  COND3X1 U12723 ( .A(n17731), .B(n16939), .C(n13788), .D(n13787), .Z(n11298)
         );
  COND1XL U12724 ( .A(Poly13[523]), .B(Poly13[396]), .C(n17298), .Z(n13790) );
  CMXI2X1 U12725 ( .A0(n18095), .A1(poly13_shifted[424]), .S(n17043), .Z(
        n13789) );
  COND4CX1 U12726 ( .A(Poly13[396]), .B(Poly13[523]), .C(n13790), .D(n13789), 
        .Z(n10650) );
  CEOXL U12727 ( .A(Poly4[50]), .B(Poly4[55]), .Z(n13791) );
  CENX1 U12728 ( .A(n16068), .B(n13791), .Z(n14484) );
  CIVX2 U12729 ( .A(n15673), .Z(n16644) );
  COND1XL U12730 ( .A(n14484), .B(Poly4[27]), .C(n16644), .Z(n13793) );
  CMXI2X1 U12731 ( .A0(n13028), .A1(Poly4[44]), .S(n12153), .Z(n13792) );
  COND4CX1 U12732 ( .A(Poly4[27]), .B(n14484), .C(n13793), .D(n13792), .Z(
        n8812) );
  CIVX2 U12733 ( .A(n15673), .Z(n17533) );
  COND1XL U12734 ( .A(Poly1[338]), .B(Poly1[200]), .C(n17533), .Z(n13795) );
  CMXI2X1 U12735 ( .A0(n18176), .A1(poly1_shifted[222]), .S(n17053), .Z(n13794) );
  COND4CX1 U12736 ( .A(Poly1[200]), .B(Poly1[338]), .C(n13795), .D(n13794), 
        .Z(n9146) );
  CENX1 U12737 ( .A(n14017), .B(n13796), .Z(n13799) );
  CIVX2 U12738 ( .A(n15673), .Z(n17215) );
  COND1XL U12739 ( .A(Poly7[410]), .B(n13799), .C(n17215), .Z(n13798) );
  CANR2X1 U12740 ( .A(n18116), .B(n17832), .C(dataselector[6]), .D(n16410), 
        .Z(n13797) );
  COND4CX1 U12741 ( .A(n13799), .B(Poly7[410]), .C(n13798), .D(n13797), .Z(
        n8789) );
  CENX1 U12742 ( .A(Poly4[53]), .B(n18214), .Z(n14112) );
  CENX1 U12743 ( .A(n13800), .B(n14614), .Z(n17580) );
  CENX1 U12744 ( .A(n14112), .B(n17580), .Z(n14493) );
  COND1XL U12745 ( .A(Poly4[25]), .B(n14493), .C(n17174), .Z(n13802) );
  CMXI2X1 U12746 ( .A0(n12013), .A1(Poly4[42]), .S(n12153), .Z(n13801) );
  COND4CX1 U12747 ( .A(n14493), .B(Poly4[25]), .C(n13802), .D(n13801), .Z(
        n8814) );
  CIVX2 U12748 ( .A(n15673), .Z(n17209) );
  COND1XL U12749 ( .A(Poly7[401]), .B(Poly7[21]), .C(n17209), .Z(n13804) );
  CMXI2X1 U12750 ( .A0(n14361), .A1(poly7_shifted[45]), .S(n12170), .Z(n13803)
         );
  COND4CX1 U12751 ( .A(Poly7[21]), .B(Poly7[401]), .C(n13804), .D(n13803), .Z(
        n10071) );
  COND1XL U12752 ( .A(Poly5[116]), .B(Poly5[121]), .C(n16985), .Z(n13806) );
  CMXI2X1 U12753 ( .A0(n12013), .A1(poly5_shifted[24]), .S(n17930), .Z(n13805)
         );
  COND4CX1 U12754 ( .A(Poly5[121]), .B(Poly5[116]), .C(n13806), .D(n13805), 
        .Z(n11516) );
  COND4CXL U12755 ( .A(Poly12[90]), .B(n14284), .C(n12013), .D(n18001), .Z(
        n13808) );
  CND2X1 U12756 ( .A(n17652), .B(poly12_shifted[122]), .Z(n13807) );
  COND3X1 U12757 ( .A(Poly12[90]), .B(n14287), .C(n13808), .D(n13807), .Z(
        n10426) );
  CMXI2X1 U12758 ( .A0(n18138), .A1(poly14_shifted[23]), .S(n18002), .Z(n13810) );
  CND2X1 U12759 ( .A(n17504), .B(Poly14[292]), .Z(n13809) );
  CND2X1 U12760 ( .A(n13810), .B(n13809), .Z(n10398) );
  CMXI2X1 U12761 ( .A0(n12010), .A1(poly8_shifted[14]), .S(n12175), .Z(n13811)
         );
  CND2X1 U12762 ( .A(n13875), .B(n13811), .Z(n11401) );
  CND2X1 U12763 ( .A(n17362), .B(Poly8[83]), .Z(n13814) );
  CMXI2X1 U12764 ( .A0(n13812), .A1(Poly8[1]), .S(n12175), .Z(n13813) );
  CND2X1 U12765 ( .A(n13814), .B(n13813), .Z(n11400) );
  COND4CX1 U12766 ( .A(Poly6[16]), .B(n13815), .C(n18095), .D(n16962), .Z(
        n13817) );
  CND2X1 U12767 ( .A(Poly6[26]), .B(n14310), .Z(n13816) );
  COND3X1 U12768 ( .A(Poly6[16]), .B(n13818), .C(n13817), .D(n13816), .Z(n9667) );
  COND1XL U12769 ( .A(Poly13[518]), .B(Poly13[273]), .C(n17620), .Z(n13820) );
  CMXI2X1 U12770 ( .A0(n14436), .A1(poly13_shifted[301]), .S(n17592), .Z(
        n13819) );
  COND4CX1 U12771 ( .A(Poly13[273]), .B(Poly13[518]), .C(n13820), .D(n13819), 
        .Z(n10773) );
  COND1XL U12772 ( .A(Poly13[515]), .B(Poly13[270]), .C(n17755), .Z(n13822) );
  COND4CX1 U12773 ( .A(Poly13[270]), .B(Poly13[515]), .C(n13822), .D(n13821), 
        .Z(n10776) );
  CMXI2XL U12774 ( .A0(n14754), .A1(poly7_shifted[18]), .S(n17564), .Z(n13824)
         );
  CND2X1 U12775 ( .A(n17655), .B(Poly7[405]), .Z(n13823) );
  CND2X1 U12776 ( .A(n13824), .B(n13823), .Z(n10098) );
  CENX1 U12777 ( .A(n16409), .B(dataselector[54]), .Z(n13825) );
  COND1XL U12778 ( .A(n13825), .B(n18228), .C(n18227), .Z(n13826) );
  CIVX1 U12779 ( .A(dataselector[61]), .Z(n16252) );
  CMXI2X1 U12780 ( .A0(n13826), .A1(n16252), .S(n16350), .Z(n8734) );
  COND1XL U12781 ( .A(Poly8[93]), .B(Poly8[78]), .C(n17998), .Z(n13828) );
  COND4CX1 U12782 ( .A(Poly8[78]), .B(Poly8[93]), .C(n13828), .D(n13827), .Z(
        n11309) );
  COND1XL U12783 ( .A(Poly8[76]), .B(Poly8[91]), .C(n17655), .Z(n13830) );
  CMXI2X1 U12784 ( .A0(n18095), .A1(Poly8[90]), .S(n17750), .Z(n13829) );
  COND4CX1 U12785 ( .A(Poly8[91]), .B(Poly8[76]), .C(n13830), .D(n13829), .Z(
        n11311) );
  COND1XL U12786 ( .A(Poly8[68]), .B(Poly8[83]), .C(n17362), .Z(n13832) );
  CMXI2X1 U12787 ( .A0(n18210), .A1(Poly8[82]), .S(n17750), .Z(n13831) );
  COND4CX1 U12788 ( .A(Poly8[83]), .B(Poly8[68]), .C(n13832), .D(n13831), .Z(
        n11319) );
  CENX1 U12789 ( .A(Poly6[19]), .B(n13833), .Z(n13836) );
  CND2X1 U12790 ( .A(n13861), .B(n13836), .Z(n13835) );
  CMXI2X1 U12791 ( .A0(n18228), .A1(Poly6[29]), .S(n14310), .Z(n13834) );
  COND3X1 U12792 ( .A(n13836), .B(n13864), .C(n13835), .D(n13834), .Z(n9664)
         );
  COND4CX1 U12793 ( .A(Poly6[29]), .B(n13861), .C(n18138), .D(n13837), .Z(
        n13839) );
  CND2X1 U12794 ( .A(n16063), .B(Poly6[39]), .Z(n13838) );
  COND3X1 U12795 ( .A(Poly6[29]), .B(n13864), .C(n13839), .D(n13838), .Z(n9654) );
  CND2X1 U12796 ( .A(n13861), .B(Poly6[11]), .Z(n13842) );
  CMXI2X1 U12797 ( .A0(n18241), .A1(Poly6[21]), .S(n13840), .Z(n13841) );
  COND3X1 U12798 ( .A(Poly6[11]), .B(n13864), .C(n13842), .D(n13841), .Z(n9672) );
  COND1XL U12799 ( .A(Poly1[340]), .B(Poly1[24]), .C(n16702), .Z(n13844) );
  CMXI2X1 U12800 ( .A0(n18053), .A1(poly1_shifted[46]), .S(n12299), .Z(n13843)
         );
  COND4CX1 U12801 ( .A(Poly1[24]), .B(Poly1[340]), .C(n13844), .D(n13843), .Z(
        n9322) );
  COND1XL U12802 ( .A(Poly12[113]), .B(Poly12[83]), .C(n16919), .Z(n13846) );
  CMXI2X1 U12803 ( .A0(poly12_shifted[115]), .A1(n18053), .S(n18001), .Z(
        n13845) );
  COND4CX1 U12804 ( .A(Poly12[83]), .B(Poly12[113]), .C(n13846), .D(n13845), 
        .Z(n10433) );
  COND1XL U12805 ( .A(Poly1[337]), .B(Poly1[199]), .C(n17238), .Z(n13848) );
  CMXI2X1 U12806 ( .A0(n18210), .A1(poly1_shifted[221]), .S(n17053), .Z(n13847) );
  COND4CX1 U12807 ( .A(Poly1[199]), .B(Poly1[337]), .C(n13848), .D(n13847), 
        .Z(n9147) );
  COND1XL U12808 ( .A(Poly1[341]), .B(Poly1[203]), .C(n16427), .Z(n13850) );
  CMXI2X1 U12809 ( .A0(n14487), .A1(poly1_shifted[225]), .S(n17053), .Z(n13849) );
  COND4CX1 U12810 ( .A(Poly1[203]), .B(Poly1[341]), .C(n13850), .D(n13849), 
        .Z(n9143) );
  COND1XL U12811 ( .A(Poly1[340]), .B(Poly1[202]), .C(n16427), .Z(n13852) );
  CMXI2X1 U12812 ( .A0(n18241), .A1(poly1_shifted[224]), .S(n17053), .Z(n13851) );
  COND4CX1 U12813 ( .A(Poly1[202]), .B(Poly1[340]), .C(n13852), .D(n13851), 
        .Z(n9144) );
  CIVX2 U12814 ( .A(n15648), .Z(n17545) );
  COND1XL U12815 ( .A(Poly0[219]), .B(Poly0[167]), .C(n17545), .Z(n13854) );
  CANR2X1 U12816 ( .A(n18249), .B(n15960), .C(poly0_shifted[203]), .D(n15671), 
        .Z(n13853) );
  COND4CX1 U12817 ( .A(Poly0[167]), .B(Poly0[219]), .C(n13854), .D(n13853), 
        .Z(n9392) );
  COND1XL U12818 ( .A(Poly5[111]), .B(Poly5[116]), .C(n17334), .Z(n13856) );
  CMXI2X1 U12819 ( .A0(n11992), .A1(poly5_shifted[19]), .S(n17930), .Z(n13855)
         );
  COND4CX1 U12820 ( .A(Poly5[116]), .B(Poly5[111]), .C(n13856), .D(n13855), 
        .Z(n11521) );
  CENX1 U12821 ( .A(Poly4[60]), .B(n18214), .Z(n15639) );
  CENX1 U12822 ( .A(Poly4[42]), .B(n15639), .Z(n13857) );
  COND1XL U12823 ( .A(Poly6[21]), .B(Poly6[49]), .C(n17072), .Z(n13860) );
  CMXI2X1 U12824 ( .A0(n12003), .A1(Poly6[31]), .S(n14310), .Z(n13859) );
  COND4CX1 U12825 ( .A(Poly6[49]), .B(Poly6[21]), .C(n13860), .D(n13859), .Z(
        n9662) );
  CND2X1 U12826 ( .A(n13861), .B(Poly6[52]), .Z(n13863) );
  CMXI2X1 U12827 ( .A0(n14754), .A1(poly6_shifted[16]), .S(n14310), .Z(n13862)
         );
  COND3X1 U12828 ( .A(Poly6[52]), .B(n13864), .C(n13863), .D(n13862), .Z(n9687) );
  CEOXL U12829 ( .A(Poly8[88]), .B(Poly8[9]), .Z(n13867) );
  COND1XL U12830 ( .A(Poly8[90]), .B(n13867), .C(n17238), .Z(n13866) );
  CMXI2X1 U12831 ( .A0(n11999), .A1(poly8_shifted[37]), .S(n12175), .Z(n13865)
         );
  COND4CX1 U12832 ( .A(n13867), .B(Poly8[90]), .C(n13866), .D(n13865), .Z(
        n11378) );
  CEOXL U12833 ( .A(Poly8[95]), .B(Poly8[14]), .Z(n13870) );
  CIVX2 U12834 ( .A(n15648), .Z(n17642) );
  COND1XL U12835 ( .A(Poly8[93]), .B(n13870), .C(n17642), .Z(n13869) );
  COND4CX1 U12836 ( .A(n13870), .B(Poly8[93]), .C(n13869), .D(n13868), .Z(
        n11373) );
  CEOX1 U12837 ( .A(Poly8[92]), .B(Poly8[11]), .Z(n13871) );
  CIVX1 U12838 ( .A(Poly8[90]), .Z(n14355) );
  CEOX1 U12839 ( .A(Poly8[3]), .B(Poly8[84]), .Z(n13876) );
  CND2X1 U12840 ( .A(n13872), .B(n13876), .Z(n13874) );
  CMXI2X1 U12841 ( .A0(n14297), .A1(poly8_shifted[31]), .S(n12175), .Z(n13873)
         );
  COND3X1 U12842 ( .A(n13876), .B(n13875), .C(n13874), .D(n13873), .Z(n11384)
         );
  CND2XL U12843 ( .A(n17298), .B(poly14_shifted[51]), .Z(n13881) );
  CND2X1 U12844 ( .A(n13878), .B(n13877), .Z(n13879) );
  CND2X1 U12845 ( .A(n17525), .B(poly14_shifted[67]), .Z(n13880) );
  COND4CX1 U12846 ( .A(n13881), .B(n17664), .C(n17525), .D(n13880), .Z(n10354)
         );
  COND1XL U12847 ( .A(n17830), .B(dataselector[29]), .C(n17535), .Z(n13884) );
  CIVDX1 U12848 ( .A(n13882), .Z0(n18252), .Z1(n15710) );
  CANR2X1 U12849 ( .A(n12004), .B(n18248), .C(n15710), .D(dataselector[36]), 
        .Z(n13883) );
  COND4CX1 U12850 ( .A(dataselector[29]), .B(n17830), .C(n13884), .D(n13883), 
        .Z(n8759) );
  CENX1 U12851 ( .A(dataselector[25]), .B(n16252), .Z(n13887) );
  COND1XL U12852 ( .A(dataselector[57]), .B(n13887), .C(n17094), .Z(n13886) );
  CANR2X1 U12853 ( .A(n18108), .B(n18248), .C(n15710), .D(dataselector[32]), 
        .Z(n13885) );
  COND4CX1 U12854 ( .A(n13887), .B(dataselector[57]), .C(n13886), .D(n13885), 
        .Z(n8763) );
  COND1XL U12855 ( .A(n17830), .B(dataselector[39]), .C(n17099), .Z(n13889) );
  CANR2X1 U12856 ( .A(n18160), .B(n18248), .C(n15710), .D(dataselector[46]), 
        .Z(n13888) );
  COND4CX1 U12857 ( .A(dataselector[39]), .B(n17830), .C(n13889), .D(n13888), 
        .Z(n8749) );
  COND1XL U12858 ( .A(Poly0[213]), .B(Poly0[16]), .C(n17705), .Z(n13891) );
  CANR2X1 U12859 ( .A(n13428), .B(n14159), .C(n17500), .D(poly0_shifted[52]), 
        .Z(n13890) );
  COND4CX1 U12860 ( .A(Poly0[16]), .B(Poly0[213]), .C(n13891), .D(n13890), .Z(
        n9543) );
  COND1XL U12861 ( .A(Poly0[217]), .B(Poly0[20]), .C(n17634), .Z(n13893) );
  CANR2X1 U12862 ( .A(n14754), .B(n14159), .C(n17500), .D(poly0_shifted[56]), 
        .Z(n13892) );
  COND4CX1 U12863 ( .A(Poly0[20]), .B(Poly0[217]), .C(n13893), .D(n13892), .Z(
        n9539) );
  COND1XL U12864 ( .A(Poly0[212]), .B(Poly0[15]), .C(n17642), .Z(n13895) );
  CANR2X1 U12865 ( .A(n14361), .B(n14159), .C(n17500), .D(poly0_shifted[51]), 
        .Z(n13894) );
  COND4CX1 U12866 ( .A(Poly0[15]), .B(Poly0[212]), .C(n13895), .D(n13894), .Z(
        n9544) );
  COND1XL U12867 ( .A(Poly0[218]), .B(Poly0[21]), .C(n17705), .Z(n13897) );
  CANR2X1 U12868 ( .A(n18138), .B(n14159), .C(n17500), .D(poly0_shifted[57]), 
        .Z(n13896) );
  COND4CX1 U12869 ( .A(Poly0[21]), .B(Poly0[218]), .C(n13897), .D(n13896), .Z(
        n9538) );
  COND1XL U12870 ( .A(Poly0[211]), .B(Poly0[14]), .C(n17466), .Z(n13899) );
  CANR2X1 U12871 ( .A(n18108), .B(n14159), .C(n17500), .D(poly0_shifted[50]), 
        .Z(n13898) );
  COND4CX1 U12872 ( .A(Poly0[14]), .B(Poly0[211]), .C(n13899), .D(n13898), .Z(
        n9545) );
  COND1XL U12873 ( .A(Poly0[215]), .B(Poly0[18]), .C(n17705), .Z(n13901) );
  CANR2X1 U12874 ( .A(n12004), .B(n14159), .C(n17500), .D(poly0_shifted[54]), 
        .Z(n13900) );
  COND4CX1 U12875 ( .A(Poly0[18]), .B(Poly0[215]), .C(n13901), .D(n13900), .Z(
        n9541) );
  COND1XL U12876 ( .A(Poly1[346]), .B(Poly1[30]), .C(n17072), .Z(n13903) );
  CMXI2X1 U12877 ( .A0(n18189), .A1(poly1_shifted[52]), .S(n12299), .Z(n13902)
         );
  COND4CX1 U12878 ( .A(Poly1[30]), .B(Poly1[346]), .C(n13903), .D(n13902), .Z(
        n9316) );
  COND1XL U12879 ( .A(Poly5[118]), .B(Poly5[83]), .C(n18047), .Z(n13906) );
  CMXI2X1 U12880 ( .A0(n14716), .A1(Poly5[97]), .S(n13904), .Z(n13905) );
  COND4CX1 U12881 ( .A(Poly5[83]), .B(Poly5[118]), .C(n13906), .D(n13905), .Z(
        n11429) );
  COND1XL U12882 ( .A(Poly5[114]), .B(Poly5[119]), .C(n16479), .Z(n13908) );
  CMXI2X1 U12883 ( .A0(n18142), .A1(poly5_shifted[22]), .S(n17930), .Z(n13907)
         );
  COND4CX1 U12884 ( .A(Poly5[119]), .B(Poly5[114]), .C(n13908), .D(n13907), 
        .Z(n11518) );
  COND1XL U12885 ( .A(Poly7[409]), .B(Poly7[29]), .C(n17288), .Z(n13910) );
  CMXI2X1 U12886 ( .A0(n18189), .A1(poly7_shifted[53]), .S(n12170), .Z(n13909)
         );
  COND4CX1 U12887 ( .A(Poly7[29]), .B(Poly7[409]), .C(n13910), .D(n13909), .Z(
        n10063) );
  COND1XL U12888 ( .A(Poly7[410]), .B(Poly7[30]), .C(n16488), .Z(n13912) );
  CMXI2X1 U12889 ( .A0(n12013), .A1(poly7_shifted[54]), .S(n12170), .Z(n13911)
         );
  COND4CX1 U12890 ( .A(Poly7[30]), .B(Poly7[410]), .C(n13912), .D(n13911), .Z(
        n10062) );
  COND1XL U12891 ( .A(Poly7[408]), .B(Poly7[28]), .C(n16323), .Z(n13914) );
  CMXI2X1 U12892 ( .A0(n18142), .A1(poly7_shifted[52]), .S(n12170), .Z(n13913)
         );
  COND4CX1 U12893 ( .A(Poly7[28]), .B(Poly7[408]), .C(n13914), .D(n13913), .Z(
        n10064) );
  COND1XL U12894 ( .A(Poly5[118]), .B(Poly5[123]), .C(n16985), .Z(n13916) );
  CMXI2X1 U12895 ( .A0(n13028), .A1(poly5_shifted[26]), .S(n17930), .Z(n13915)
         );
  COND4CX1 U12896 ( .A(Poly5[123]), .B(Poly5[118]), .C(n13916), .D(n13915), 
        .Z(n11514) );
  COND1XL U12897 ( .A(Poly7[48]), .B(Poly7[399]), .C(n17094), .Z(n13918) );
  COND4CX1 U12898 ( .A(Poly7[399]), .B(Poly7[48]), .C(n13918), .D(n13917), .Z(
        n10044) );
  COND1XL U12899 ( .A(Poly5[115]), .B(Poly5[120]), .C(n16488), .Z(n13920) );
  CMXI2X1 U12900 ( .A0(n18189), .A1(poly5_shifted[23]), .S(n17932), .Z(n13919)
         );
  COND4CX1 U12901 ( .A(Poly5[120]), .B(Poly5[115]), .C(n13920), .D(n13919), 
        .Z(n11517) );
  COND1XL U12902 ( .A(\dataselector_shifted[0] ), .B(Poly7[24]), .C(n17121), 
        .Z(n13922) );
  CMXI2X1 U12903 ( .A0(n12004), .A1(poly7_shifted[48]), .S(n12170), .Z(n13921)
         );
  COND4CX1 U12904 ( .A(Poly7[24]), .B(\dataselector_shifted[0] ), .C(n13922), 
        .D(n13921), .Z(n10068) );
  COND1XL U12905 ( .A(Poly7[402]), .B(Poly7[51]), .C(n17280), .Z(n13924) );
  CMXI2X1 U12906 ( .A0(n14436), .A1(poly7_shifted[75]), .S(n12170), .Z(n13923)
         );
  COND4CX1 U12907 ( .A(Poly7[51]), .B(Poly7[402]), .C(n13924), .D(n13923), .Z(
        n10041) );
  COND1XL U12908 ( .A(Poly7[406]), .B(Poly7[26]), .C(n17198), .Z(n13926) );
  CMXI2X1 U12909 ( .A0(n14754), .A1(poly7_shifted[50]), .S(n12170), .Z(n13925)
         );
  COND4CX1 U12910 ( .A(Poly7[26]), .B(Poly7[406]), .C(n13926), .D(n13925), .Z(
        n10066) );
  CENX1 U12911 ( .A(n14615), .B(n13927), .Z(n14620) );
  CENX1 U12912 ( .A(n15651), .B(n13928), .Z(n13929) );
  CENX1 U12913 ( .A(n14620), .B(n13929), .Z(n15865) );
  COND1XL U12914 ( .A(Poly4[16]), .B(n15865), .C(n17290), .Z(n13931) );
  CMXI2X1 U12915 ( .A0(n14765), .A1(Poly4[33]), .S(n12153), .Z(n13930) );
  COND4CX1 U12916 ( .A(n15865), .B(Poly4[16]), .C(n13931), .D(n13930), .Z(
        n8823) );
  COND1XL U12917 ( .A(Poly7[25]), .B(Poly7[405]), .C(n16488), .Z(n13933) );
  CMXI2X1 U12918 ( .A0(n11982), .A1(poly7_shifted[49]), .S(n12170), .Z(n13932)
         );
  COND4CX1 U12919 ( .A(Poly7[405]), .B(Poly7[25]), .C(n13933), .D(n13932), .Z(
        n10067) );
  CIVX2 U12920 ( .A(n15673), .Z(n17178) );
  COND1XL U12921 ( .A(Poly7[407]), .B(Poly7[27]), .C(n17178), .Z(n13935) );
  CMXI2X1 U12922 ( .A0(n18138), .A1(poly7_shifted[51]), .S(n12170), .Z(n13934)
         );
  COND4CX1 U12923 ( .A(Poly7[27]), .B(Poly7[407]), .C(n13935), .D(n13934), .Z(
        n10065) );
  COND1XL U12924 ( .A(dataselector[38]), .B(n14022), .C(n17535), .Z(n13937) );
  CANR2X1 U12925 ( .A(n18219), .B(n18248), .C(n16350), .D(dataselector[45]), 
        .Z(n13936) );
  COND4CX1 U12926 ( .A(n14022), .B(dataselector[38]), .C(n13937), .D(n13936), 
        .Z(n8750) );
  CENX1 U12927 ( .A(n16385), .B(n14943), .Z(n13991) );
  COND1XL U12928 ( .A(n13991), .B(dataselector[36]), .C(n17063), .Z(n13939) );
  CANR2X1 U12929 ( .A(n16381), .B(n18248), .C(n16350), .D(dataselector[43]), 
        .Z(n13938) );
  COND4CX1 U12930 ( .A(dataselector[36]), .B(n13991), .C(n13939), .D(n13938), 
        .Z(n8752) );
  CMXI2X1 U12931 ( .A0(n18053), .A1(poly15_shifted[50]), .S(n17376), .Z(n13944) );
  CIVX2 U12932 ( .A(n18040), .Z(n16796) );
  CIVX2 U12933 ( .A(n13940), .Z(n18042) );
  CENX1 U12934 ( .A(Poly15[52]), .B(Poly15[53]), .Z(n13941) );
  CENX1 U12935 ( .A(Poly15[20]), .B(n13941), .Z(n13942) );
  CMXI2X1 U12936 ( .A0(n16796), .A1(n18042), .S(n13942), .Z(n13943) );
  CND2X1 U12937 ( .A(n13944), .B(n13943), .Z(n9602) );
  CIVX2 U12938 ( .A(n17259), .Z(n17348) );
  CND2X1 U12939 ( .A(n14848), .B(entrophy[18]), .Z(n14965) );
  CND2X1 U12940 ( .A(n17759), .B(entrophy[22]), .Z(n14683) );
  CNR2X2 U12941 ( .A(n14226), .B(n13947), .Z(n14982) );
  CND2X1 U12942 ( .A(n15206), .B(datain[4]), .Z(n14416) );
  CNR2X1 U12943 ( .A(n15218), .B(n14453), .Z(n14962) );
  CIVX1 U12944 ( .A(n14962), .Z(n13950) );
  CND2X1 U12945 ( .A(n14998), .B(n13950), .Z(n13952) );
  CAN2XL U12946 ( .A(n13945), .B(entrophy[2]), .Z(n13951) );
  CND3XL U12947 ( .A(n15274), .B(n17804), .C(entrophy[31]), .Z(n13975) );
  CND2XL U12948 ( .A(n17829), .B(scrambler[5]), .Z(n13955) );
  CND2XL U12949 ( .A(n15334), .B(n13955), .Z(n13967) );
  CNR2X1 U12950 ( .A(n15168), .B(n14999), .Z(n13957) );
  CIVXL U12951 ( .A(n13955), .Z(n13956) );
  CANR3X1 U12952 ( .A(n15130), .B(dataselector[14]), .C(n13957), .D(n13956), 
        .Z(n13960) );
  CIVDX1 U12953 ( .A(n13958), .Z0(n17776), .Z1(n14559) );
  COR2X1 U12954 ( .A(n15219), .B(n14559), .Z(n14705) );
  CNR2X1 U12955 ( .A(n14969), .B(n14686), .Z(n14838) );
  CND2X1 U12956 ( .A(n15206), .B(dataselector[14]), .Z(n15075) );
  CNR2XL U12957 ( .A(n15075), .B(n14659), .Z(n13959) );
  CND2XL U12958 ( .A(n17804), .B(entrophy[13]), .Z(n14930) );
  CIVX1 U12959 ( .A(n14976), .Z(n15104) );
  CIVX1 U12960 ( .A(datain[6]), .Z(n14471) );
  CNR2X1 U12961 ( .A(n15149), .B(n14471), .Z(n13963) );
  CND2X1 U12962 ( .A(n14826), .B(entrophy[8]), .Z(n14689) );
  CIVX1 U12963 ( .A(n14689), .Z(n13961) );
  CIVX2 U12964 ( .A(n15327), .Z(n14917) );
  COND11X1 U12965 ( .A(n13963), .B(n13962), .C(n13961), .D(n14917), .Z(n13964)
         );
  COND1XL U12966 ( .A(n14930), .B(n15104), .C(n13964), .Z(n13965) );
  CANR1X1 U12967 ( .A(n13967), .B(n13966), .C(n13965), .Z(n13974) );
  CNR2X1 U12968 ( .A(n15351), .B(n14850), .Z(n15018) );
  CIVXL U12969 ( .A(n15018), .Z(n13968) );
  CND2XL U12970 ( .A(n15256), .B(entrophy[26]), .Z(n15120) );
  CNR2X1 U12971 ( .A(n15218), .B(n14886), .Z(n14474) );
  CIVX1 U12972 ( .A(n14474), .Z(n15053) );
  CND3XL U12973 ( .A(n13968), .B(n15120), .C(n15053), .Z(n13972) );
  CIVX1 U12974 ( .A(n13969), .Z(n13970) );
  CIVDX1 U12975 ( .A(n15200), .Z0(n12520), .Z1(n14857) );
  CND2X1 U12976 ( .A(n14857), .B(entrophy[28]), .Z(n14068) );
  CND2X1 U12977 ( .A(n12019), .B(datain[2]), .Z(n17779) );
  CND3XL U12978 ( .A(n13970), .B(n14068), .C(n17779), .Z(n13971) );
  CND2X1 U12979 ( .A(n15035), .B(entrophy[25]), .Z(n15124) );
  CNR2X1 U12980 ( .A(n15124), .B(n14085), .Z(n14957) );
  COND11X1 U12981 ( .A(n13972), .B(n13971), .C(n14957), .D(n15145), .Z(n13973)
         );
  CND4X1 U12982 ( .A(n13976), .B(n13975), .C(n13974), .D(n13973), .Z(n8705) );
  CIVXL U12983 ( .A(n16274), .Z(n13979) );
  CND2X1 U12984 ( .A(n15880), .B(Poly0[109]), .Z(n13978) );
  CND2X1 U12985 ( .A(n17598), .B(poly0_shifted[109]), .Z(n13977) );
  COND3X1 U12986 ( .A(n13979), .B(n17090), .C(n13978), .D(n13977), .Z(n9468)
         );
  CND2X1 U12987 ( .A(n12997), .B(poly12_shifted[29]), .Z(n13981) );
  CND2XL U12988 ( .A(n17504), .B(Poly12[124]), .Z(n13980) );
  COND3X1 U12989 ( .A(n12997), .B(n17090), .C(n13981), .D(n13980), .Z(n10519)
         );
  COND1XL U12990 ( .A(Poly13[526]), .B(Poly13[281]), .C(n18234), .Z(n13983) );
  CMXI2X1 U12991 ( .A0(n18138), .A1(poly13_shifted[309]), .S(n17615), .Z(
        n13982) );
  COND4CX1 U12992 ( .A(Poly13[281]), .B(Poly13[526]), .C(n13983), .D(n13982), 
        .Z(n10765) );
  COND1XL U12993 ( .A(Poly13[522]), .B(Poly13[277]), .C(n16919), .Z(n13985) );
  CMXI2X1 U12994 ( .A0(n18053), .A1(poly13_shifted[305]), .S(n17615), .Z(
        n13984) );
  COND4CX1 U12995 ( .A(Poly13[277]), .B(Poly13[522]), .C(n13985), .D(n13984), 
        .Z(n10769) );
  CIVXL U12996 ( .A(Poly13[527]), .Z(n13986) );
  CND2X1 U12997 ( .A(n12997), .B(poly12_shifted[21]), .Z(n13988) );
  CND2XL U12998 ( .A(n17755), .B(Poly12[116]), .Z(n13987) );
  COND3X1 U12999 ( .A(n12997), .B(n11985), .C(n13988), .D(n13987), .Z(n10527)
         );
  COND1XL U13000 ( .A(dataselector[20]), .B(n13991), .C(n17094), .Z(n13990) );
  CANR2X1 U13001 ( .A(n18099), .B(n17832), .C(dataselector[27]), .D(n16410), 
        .Z(n13989) );
  COND4CX1 U13002 ( .A(n13991), .B(dataselector[20]), .C(n13990), .D(n13989), 
        .Z(n8768) );
  COND1XL U13003 ( .A(dataselector[16]), .B(n15919), .C(n17535), .Z(n13993) );
  CANR2X1 U13004 ( .A(n11999), .B(n17832), .C(dataselector[23]), .D(n16410), 
        .Z(n13992) );
  COND4CX1 U13005 ( .A(n15919), .B(dataselector[16]), .C(n13993), .D(n13992), 
        .Z(n8772) );
  COND1XL U13006 ( .A(dataselector[17]), .B(n17828), .C(n17535), .Z(n13996) );
  CANR2X1 U13007 ( .A(n13994), .B(n17832), .C(dataselector[24]), .D(n16410), 
        .Z(n13995) );
  COND4CX1 U13008 ( .A(n17828), .B(dataselector[17]), .C(n13996), .D(n13995), 
        .Z(n8771) );
  CND2X1 U13009 ( .A(n14005), .B(Poly6[33]), .Z(n13998) );
  CMXI2X1 U13010 ( .A0(n16381), .A1(Poly6[43]), .S(n14166), .Z(n13997) );
  COND3X1 U13011 ( .A(Poly6[33]), .B(n14008), .C(n13998), .D(n13997), .Z(n9650) );
  CND2X1 U13012 ( .A(n14005), .B(Poly6[46]), .Z(n14000) );
  CMXI2X1 U13013 ( .A0(n11988), .A1(poly6_shifted[15]), .S(n14310), .Z(n13999)
         );
  COND3X1 U13014 ( .A(Poly6[46]), .B(n14008), .C(n14000), .D(n13999), .Z(n9688) );
  COND4CX1 U13015 ( .A(Poly6[15]), .B(n14005), .C(n17934), .D(n16962), .Z(
        n14002) );
  CND2X1 U13016 ( .A(Poly6[25]), .B(n14310), .Z(n14001) );
  COND3X1 U13017 ( .A(Poly6[15]), .B(n14008), .C(n14002), .D(n14001), .Z(n9668) );
  COND4CXL U13018 ( .A(Poly6[0]), .B(n14005), .C(n12013), .D(n16962), .Z(
        n14004) );
  CND2X1 U13019 ( .A(n14310), .B(Poly6[10]), .Z(n14003) );
  COND3X1 U13020 ( .A(Poly6[0]), .B(n14008), .C(n14004), .D(n14003), .Z(n9683)
         );
  CND2X1 U13021 ( .A(n14005), .B(Poly6[23]), .Z(n14007) );
  CMXI2X1 U13022 ( .A0(n14361), .A1(Poly6[33]), .S(n14166), .Z(n14006) );
  COND3X1 U13023 ( .A(Poly6[23]), .B(n14008), .C(n14007), .D(n14006), .Z(n9660) );
  CND2X1 U13024 ( .A(n18082), .B(n17832), .Z(n14011) );
  CEOXL U13025 ( .A(dataselector[13]), .B(dataselector[59]), .Z(n14009) );
  CANR2X1 U13026 ( .A(n16410), .B(dataselector[20]), .C(n17533), .D(n14009), 
        .Z(n14010) );
  CND2X1 U13027 ( .A(n14011), .B(n14010), .Z(n8775) );
  COND1XL U13028 ( .A(n14014), .B(Poly11[56]), .C(n17508), .Z(n14013) );
  CMXI2X1 U13029 ( .A0(n18138), .A1(Poly11[71]), .S(n15843), .Z(n14012) );
  COND4CX1 U13030 ( .A(Poly11[56]), .B(n14014), .C(n14013), .D(n14012), .Z(
        n11118) );
  COND1XL U13031 ( .A(Poly12[114]), .B(Poly12[18]), .C(n17266), .Z(n14016) );
  CMXI2X1 U13032 ( .A0(n13428), .A1(Poly12[34]), .S(n12598), .Z(n14015) );
  COND4CX1 U13033 ( .A(Poly12[18]), .B(Poly12[114]), .C(n14016), .D(n14015), 
        .Z(n10498) );
  CEOX1 U13034 ( .A(n14017), .B(dataselector[63]), .Z(n18247) );
  COND1XL U13035 ( .A(Poly7[408]), .B(n18247), .C(n17105), .Z(n14019) );
  CANR2X1 U13036 ( .A(n12004), .B(n17832), .C(dataselector[4]), .D(n16410), 
        .Z(n14018) );
  COND4CX1 U13037 ( .A(n18247), .B(Poly7[408]), .C(n14019), .D(n14018), .Z(
        n8791) );
  COND1XL U13038 ( .A(n14022), .B(dataselector[22]), .C(n17063), .Z(n14021) );
  CANR2X1 U13039 ( .A(n18228), .B(n17832), .C(dataselector[29]), .D(n16410), 
        .Z(n14020) );
  COND4CX1 U13040 ( .A(dataselector[22]), .B(n14022), .C(n14021), .D(n14020), 
        .Z(n8766) );
  COND1XL U13041 ( .A(dataselector[61]), .B(dataselector[15]), .C(n17535), .Z(
        n14024) );
  CANR2X1 U13042 ( .A(n18034), .B(n17832), .C(dataselector[22]), .D(n16410), 
        .Z(n14023) );
  COND4CX1 U13043 ( .A(dataselector[15]), .B(dataselector[61]), .C(n14024), 
        .D(n14023), .Z(n8773) );
  CND2X1 U13044 ( .A(n15256), .B(entrophy[6]), .Z(n15267) );
  CND2X1 U13045 ( .A(n14695), .B(entrophy[8]), .Z(n14374) );
  CND3XL U13046 ( .A(n14965), .B(n15267), .C(n14374), .Z(n14027) );
  CND2X1 U13047 ( .A(n15319), .B(datain[7]), .Z(n14600) );
  COND3X1 U13048 ( .A(n15351), .B(n14926), .C(n14600), .D(n14025), .Z(n14026)
         );
  CANR3X1 U13049 ( .A(n15119), .B(entrophy[30]), .C(n14027), .D(n14026), .Z(
        n14045) );
  CIVX1 U13050 ( .A(n14093), .Z(n14030) );
  CND2X1 U13051 ( .A(n14857), .B(entrophy[0]), .Z(n14582) );
  CND2X1 U13052 ( .A(n17759), .B(entrophy[10]), .Z(n14847) );
  CIVX2 U13053 ( .A(entrophy[17]), .Z(n15229) );
  CNR2X1 U13054 ( .A(n15351), .B(n15229), .Z(n14130) );
  CIVX1 U13055 ( .A(n14130), .Z(n14029) );
  CND2X1 U13056 ( .A(n12019), .B(datain[7]), .Z(n15060) );
  CIVX1 U13057 ( .A(dataselector[25]), .Z(n15798) );
  CND2X1 U13058 ( .A(n17768), .B(n15798), .Z(n15191) );
  CND8X1 U13059 ( .A(n14030), .B(n14582), .C(n14847), .D(n14029), .E(n15060), 
        .F(n15191), .G(n14028), .H(n14075), .Z(n14037) );
  CNR2X1 U13060 ( .A(n14969), .B(n14659), .Z(n15099) );
  CIVXL U13061 ( .A(n15099), .Z(n14031) );
  CND2X1 U13062 ( .A(n14695), .B(entrophy[18]), .Z(n17766) );
  CND2X1 U13063 ( .A(n15256), .B(entrophy[0]), .Z(n14902) );
  CAN4X1 U13064 ( .A(n14031), .B(n17766), .C(n14902), .D(n14824), .Z(n14035)
         );
  CND2X1 U13065 ( .A(n15319), .B(entrophy[8]), .Z(n14638) );
  COR2XL U13066 ( .A(n14472), .B(n15352), .Z(n14032) );
  CND2X1 U13067 ( .A(n14638), .B(n14032), .Z(n15203) );
  CIVX1 U13068 ( .A(n15203), .Z(n14034) );
  CND2X1 U13069 ( .A(n14033), .B(datain[3]), .Z(n14229) );
  CND2X1 U13070 ( .A(n14084), .B(entrophy[3]), .Z(n15171) );
  CND4X1 U13071 ( .A(n14035), .B(n14034), .C(n14229), .D(n15171), .Z(n14036)
         );
  CANR2X1 U13072 ( .A(n15145), .B(n14037), .C(n12216), .D(n14036), .Z(n14044)
         );
  CIVX1 U13073 ( .A(n15071), .Z(n14039) );
  CND2X1 U13074 ( .A(n15206), .B(entrophy[26]), .Z(n15025) );
  CIVXL U13075 ( .A(n15025), .Z(n14038) );
  CNR2X1 U13076 ( .A(n14969), .B(n14465), .Z(n14091) );
  CNR4X1 U13077 ( .A(n14039), .B(n14038), .C(n15193), .D(n14091), .Z(n14041)
         );
  CANR1XL U13078 ( .A(entrophy[14]), .B(n14131), .C(n15005), .Z(n14040) );
  CND2X1 U13079 ( .A(n14857), .B(entrophy[16]), .Z(n14802) );
  CND4X1 U13080 ( .A(n14041), .B(n14040), .C(n14600), .D(n14802), .Z(n14042)
         );
  CANR2XL U13081 ( .A(n14042), .B(n15220), .C(scrambler[31]), .D(n17744), .Z(
        n14043) );
  COND3X1 U13082 ( .A(n14045), .B(n15236), .C(n14044), .D(n14043), .Z(n8731)
         );
  CENX1 U13083 ( .A(Poly15[51]), .B(Poly15[52]), .Z(n14046) );
  CENX1 U13084 ( .A(Poly15[19]), .B(n14046), .Z(n14049) );
  COND1XL U13085 ( .A(Poly15[45]), .B(n14049), .C(n17094), .Z(n14048) );
  CMXI2X1 U13086 ( .A0(n12415), .A1(poly15_shifted[49]), .S(n17376), .Z(n14047) );
  COND4CX1 U13087 ( .A(n14049), .B(Poly15[45]), .C(n14048), .D(n14047), .Z(
        n9603) );
  COND1XL U13088 ( .A(Poly1[343]), .B(Poly1[158]), .C(n17613), .Z(n14051) );
  CMXI2X1 U13089 ( .A0(n12001), .A1(poly1_shifted[180]), .S(n12210), .Z(n14050) );
  COND4CX1 U13090 ( .A(Poly1[158]), .B(Poly1[343]), .C(n14051), .D(n14050), 
        .Z(n9188) );
  COND1XL U13091 ( .A(Poly1[337]), .B(Poly1[152]), .C(n17545), .Z(n14053) );
  CMXI2X1 U13092 ( .A0(n18053), .A1(poly1_shifted[174]), .S(n12210), .Z(n14052) );
  COND4CX1 U13093 ( .A(Poly1[152]), .B(Poly1[337]), .C(n14053), .D(n14052), 
        .Z(n9194) );
  COND1XL U13094 ( .A(Poly1[344]), .B(Poly1[159]), .C(n17560), .Z(n14055) );
  CMXI2X1 U13095 ( .A0(n12013), .A1(poly1_shifted[181]), .S(n12210), .Z(n14054) );
  COND4CX1 U13096 ( .A(Poly1[159]), .B(Poly1[344]), .C(n14055), .D(n14054), 
        .Z(n9187) );
  COND1XL U13097 ( .A(Poly1[346]), .B(Poly1[161]), .C(n17072), .Z(n14057) );
  CMXI2X1 U13098 ( .A0(n13028), .A1(poly1_shifted[183]), .S(n12210), .Z(n14056) );
  COND4CX1 U13099 ( .A(Poly1[161]), .B(Poly1[346]), .C(n14057), .D(n14056), 
        .Z(n9185) );
  COND1XL U13100 ( .A(Poly1[336]), .B(Poly1[151]), .C(n16372), .Z(n14059) );
  CMXI2X1 U13101 ( .A0(n12415), .A1(poly1_shifted[173]), .S(n12210), .Z(n14058) );
  COND4CX1 U13102 ( .A(Poly1[151]), .B(Poly1[336]), .C(n14059), .D(n14058), 
        .Z(n9195) );
  COND1XL U13103 ( .A(Poly1[345]), .B(Poly1[160]), .C(n18047), .Z(n14061) );
  CMXI2X1 U13104 ( .A0(n16381), .A1(poly1_shifted[182]), .S(n12210), .Z(n14060) );
  COND4CX1 U13105 ( .A(Poly1[160]), .B(Poly1[345]), .C(n14061), .D(n14060), 
        .Z(n9186) );
  COND1XL U13106 ( .A(Poly1[338]), .B(Poly1[153]), .C(n17449), .Z(n14063) );
  CMXI2X1 U13107 ( .A0(n12004), .A1(poly1_shifted[175]), .S(n12210), .Z(n14062) );
  COND4CX1 U13108 ( .A(Poly1[153]), .B(Poly1[338]), .C(n14063), .D(n14062), 
        .Z(n9193) );
  COND1XL U13109 ( .A(Poly9[105]), .B(Poly9[84]), .C(n17280), .Z(n14065) );
  CMXI2X1 U13110 ( .A0(n14436), .A1(poly9_shifted[106]), .S(n17955), .Z(n14064) );
  COND4CX1 U13111 ( .A(Poly9[84]), .B(Poly9[105]), .C(n14065), .D(n14064), .Z(
        n11210) );
  CMXI2X1 U13112 ( .A0(n18142), .A1(poly4_shifted[25]), .S(n18230), .Z(n14067)
         );
  CND2X1 U13113 ( .A(n17094), .B(n14614), .Z(n14066) );
  CND2X1 U13114 ( .A(n14067), .B(n14066), .Z(n8848) );
  CND3XL U13115 ( .A(n14880), .B(n18234), .C(entrophy[26]), .Z(n17773) );
  CIVX2 U13116 ( .A(n14068), .Z(n14069) );
  CNR2X1 U13117 ( .A(n15334), .B(n14788), .Z(n15047) );
  COND1X1 U13118 ( .A(n14950), .B(n14069), .C(n15047), .Z(n14072) );
  CND4X1 U13119 ( .A(n14070), .B(n14670), .C(n15309), .D(n11969), .Z(n14071)
         );
  COND3X1 U13120 ( .A(n15334), .B(n17773), .C(n14072), .D(n14071), .Z(n14077)
         );
  CNR2X1 U13121 ( .A(n15283), .B(n15219), .Z(n14372) );
  CIVX2 U13122 ( .A(n14073), .Z(n14214) );
  COND1XL U13123 ( .A(n14372), .B(n14214), .C(n12216), .Z(n14074) );
  CND2X1 U13124 ( .A(n17797), .B(entrophy[29]), .Z(n14643) );
  CIVX2 U13125 ( .A(n14643), .Z(n14576) );
  CND2X1 U13126 ( .A(n14576), .B(n14672), .Z(n15009) );
  CND2X1 U13127 ( .A(n17759), .B(entrophy[25]), .Z(n14414) );
  CIVXL U13128 ( .A(n14372), .Z(n14079) );
  CAN4X1 U13129 ( .A(n15009), .B(n14414), .C(n14080), .D(n14079), .Z(n14082)
         );
  CND2X1 U13130 ( .A(n15319), .B(entrophy[12]), .Z(n15095) );
  CAN4X1 U13131 ( .A(n14082), .B(n14081), .C(n14397), .D(n15095), .Z(n14083)
         );
  CNR2X1 U13132 ( .A(n14083), .B(n17763), .Z(n14099) );
  CND2X1 U13133 ( .A(n14084), .B(entrophy[1]), .Z(n14570) );
  CNR2X1 U13134 ( .A(n15334), .B(n17784), .Z(n15033) );
  CANR2X1 U13135 ( .A(n17770), .B(n15033), .C(n15309), .D(n15205), .Z(n14087)
         );
  CNR2IX2 U13136 ( .B(n14652), .A(n11969), .Z(n17767) );
  CAN2X1 U13137 ( .A(n17767), .B(n14085), .Z(n15034) );
  CNR2X1 U13138 ( .A(n15334), .B(n15229), .Z(n14951) );
  COND3X1 U13139 ( .A(n14570), .B(n17785), .C(n14087), .D(n14086), .Z(n14088)
         );
  CIVX2 U13140 ( .A(n14088), .Z(n14097) );
  CNR2X2 U13141 ( .A(n15351), .B(n14908), .Z(n14574) );
  COND4CXL U13142 ( .A(entrophy[28]), .B(n17759), .C(n14574), .D(n15309), .Z(
        n14089) );
  COND11XL U13143 ( .A(n17785), .B(n14230), .C(n14795), .D(n14089), .Z(n14090)
         );
  CIVX2 U13144 ( .A(n14090), .Z(n14096) );
  CND2X1 U13145 ( .A(n14084), .B(entrophy[30]), .Z(n14988) );
  CIVX1 U13146 ( .A(n14988), .Z(n14094) );
  CND2X1 U13147 ( .A(n17620), .B(entrophy[21]), .Z(n14968) );
  COND11X1 U13148 ( .A(n14094), .B(n14093), .C(n14092), .D(n14917), .Z(n14095)
         );
  CND3XL U13149 ( .A(n14097), .B(n14096), .C(n14095), .Z(n14098) );
  CNR2X1 U13150 ( .A(n14099), .B(n14098), .Z(n14100) );
  CND2X1 U13151 ( .A(n14101), .B(n14100), .Z(n8702) );
  COND1XL U13152 ( .A(Poly13[516]), .B(Poly13[157]), .C(n17362), .Z(n14103) );
  CMXI2X1 U13153 ( .A0(n16381), .A1(poly13_shifted[185]), .S(n13014), .Z(
        n14102) );
  COND4CX1 U13154 ( .A(Poly13[157]), .B(Poly13[516]), .C(n14103), .D(n14102), 
        .Z(n10889) );
  CEOX1 U13155 ( .A(Poly12[29]), .B(Poly12[125]), .Z(n14106) );
  CND2X1 U13156 ( .A(n14107), .B(n14106), .Z(n14105) );
  CMXI2X1 U13157 ( .A0(n18219), .A1(poly12_shifted[61]), .S(n12598), .Z(n14104) );
  COND3X1 U13158 ( .A(n14106), .B(n14110), .C(n14105), .D(n14104), .Z(n10487)
         );
  CEOX1 U13159 ( .A(Poly12[111]), .B(Poly12[22]), .Z(n14111) );
  CND2X1 U13160 ( .A(n14107), .B(n14111), .Z(n14109) );
  CMXI2X1 U13161 ( .A0(n18116), .A1(poly12_shifted[54]), .S(n12598), .Z(n14108) );
  COND3X1 U13162 ( .A(n14111), .B(n14110), .C(n14109), .D(n14108), .Z(n10494)
         );
  CMXI2X1 U13163 ( .A0(n12001), .A1(poly4_shifted[26]), .S(n18230), .Z(n14114)
         );
  CAN2X1 U13164 ( .A(n16947), .B(Poly4[57]), .Z(n18220) );
  CNR2X1 U13165 ( .A(n17495), .B(Poly4[57]), .Z(n18221) );
  CMXI2X1 U13166 ( .A0(n18220), .A1(n18221), .S(n14112), .Z(n14113) );
  CND2X1 U13167 ( .A(n14114), .B(n14113), .Z(n8847) );
  CMXI2X1 U13168 ( .A0(n18206), .A1(poly4_shifted[32]), .S(n18230), .Z(n14115)
         );
  CND2X1 U13169 ( .A(n17285), .B(Poly4[59]), .Z(n18218) );
  CND2X1 U13170 ( .A(n14115), .B(n18218), .Z(n8841) );
  COND1XL U13171 ( .A(Poly13[514]), .B(Poly13[155]), .C(n17508), .Z(n14117) );
  CMXI2X1 U13172 ( .A0(n18189), .A1(poly13_shifted[183]), .S(n13014), .Z(
        n14116) );
  COND4CX1 U13173 ( .A(Poly13[155]), .B(Poly13[514]), .C(n14117), .D(n14116), 
        .Z(n10891) );
  CND2X1 U13174 ( .A(n17930), .B(poly5_shifted[37]), .Z(n14119) );
  CND2XL U13175 ( .A(n17458), .B(poly5_shifted[23]), .Z(n14118) );
  COND3X1 U13176 ( .A(n17930), .B(n12000), .C(n14119), .D(n14118), .Z(n11503)
         );
  COND1XL U13177 ( .A(Poly13[520]), .B(Poly13[161]), .C(n17538), .Z(n14121) );
  CMXI2X1 U13178 ( .A0(n18206), .A1(poly13_shifted[189]), .S(n13014), .Z(
        n14120) );
  COND4CX1 U13179 ( .A(Poly13[161]), .B(Poly13[520]), .C(n14121), .D(n14120), 
        .Z(n10885) );
  CMXI2X1 U13180 ( .A0(n14361), .A1(poly14_shifted[17]), .S(n18002), .Z(n14123) );
  CND2X1 U13181 ( .A(n17266), .B(Poly14[286]), .Z(n14122) );
  CND2X1 U13182 ( .A(n14123), .B(n14122), .Z(n10404) );
  CMXI2X1 U13183 ( .A0(n11992), .A1(poly14_shifted[21]), .S(n18002), .Z(n14125) );
  CND2X1 U13184 ( .A(n17466), .B(Poly14[290]), .Z(n14124) );
  CND2X1 U13185 ( .A(n14125), .B(n14124), .Z(n10400) );
  CMXI2X1 U13186 ( .A0(n18142), .A1(poly14_shifted[24]), .S(n18002), .Z(n14127) );
  CND2X1 U13187 ( .A(n17383), .B(Poly14[293]), .Z(n14126) );
  CND2X1 U13188 ( .A(n14127), .B(n14126), .Z(n10397) );
  CND2X1 U13189 ( .A(n17759), .B(entrophy[8]), .Z(n15142) );
  CND2X1 U13190 ( .A(n15256), .B(entrophy[19]), .Z(n14417) );
  CIVXL U13191 ( .A(n15195), .Z(n14128) );
  CND2X1 U13192 ( .A(n17776), .B(entrophy[9]), .Z(n14905) );
  CND2X1 U13193 ( .A(n12019), .B(datain[6]), .Z(n15141) );
  CAN8X1 U13194 ( .A(n15142), .B(n14417), .C(n14128), .D(n15115), .E(n15063), 
        .F(n14905), .G(n15141), .H(n15114), .Z(n14147) );
  CNR2X1 U13195 ( .A(n15283), .B(n14968), .Z(n15022) );
  COR4X1 U13196 ( .A(n14866), .B(n15022), .C(n14130), .D(n14129), .Z(n14138)
         );
  CIVX1 U13197 ( .A(n14593), .Z(n14895) );
  CND2X1 U13198 ( .A(n14131), .B(entrophy[18]), .Z(n14375) );
  CND2X1 U13199 ( .A(n14857), .B(entrophy[19]), .Z(n14837) );
  COND3X1 U13200 ( .A(n14895), .B(n15211), .C(n14375), .D(n14837), .Z(n14137)
         );
  CND2X1 U13201 ( .A(n17759), .B(datain[4]), .Z(n14589) );
  COND1XL U13202 ( .A(n14561), .B(n12459), .C(n14589), .Z(n15284) );
  CNR2X1 U13203 ( .A(n14559), .B(n14999), .Z(n15006) );
  CNR2XL U13204 ( .A(n14226), .B(n14808), .Z(n14135) );
  CIVX2 U13205 ( .A(n14416), .Z(n14409) );
  CNR2X1 U13206 ( .A(n14546), .B(n14133), .Z(n14575) );
  COR8X1 U13207 ( .A(n15284), .B(n14652), .C(n15006), .D(n14135), .E(n14409), 
        .F(n14962), .G(n14134), .H(n14575), .Z(n14136) );
  COND3X1 U13208 ( .A(n14138), .B(n14137), .C(n14136), .D(n14875), .Z(n14146)
         );
  CIVX2 U13209 ( .A(n14913), .Z(n14538) );
  CNR3X1 U13210 ( .A(n14538), .B(n14139), .C(n15301), .Z(n15059) );
  CIVX2 U13211 ( .A(entrophy[29]), .Z(n14927) );
  CNR2X1 U13212 ( .A(n15283), .B(n14927), .Z(n15313) );
  CND2X1 U13213 ( .A(n15297), .B(n15150), .Z(n14707) );
  CND4XL U13214 ( .A(n14998), .B(n14140), .C(n15095), .D(n14375), .Z(n14141)
         );
  COR4X1 U13215 ( .A(n15059), .B(n15313), .C(n14707), .D(n14141), .Z(n14144)
         );
  CND2XL U13216 ( .A(n17744), .B(scrambler[6]), .Z(n14142) );
  COND11X1 U13217 ( .A(n14886), .B(n14977), .C(n14935), .D(n14142), .Z(n14143)
         );
  COND3X1 U13218 ( .A(n14147), .B(n12055), .C(n14146), .D(n14145), .Z(n8706)
         );
  COND1XL U13219 ( .A(Poly5[123]), .B(Poly5[88]), .C(n17094), .Z(n14149) );
  CMXI2X1 U13220 ( .A0(n14754), .A1(Poly5[102]), .S(n12016), .Z(n14148) );
  COND4CX1 U13221 ( .A(Poly5[88]), .B(Poly5[123]), .C(n14149), .D(n14148), .Z(
        n11424) );
  COND1XL U13222 ( .A(Poly1[340]), .B(Poly1[155]), .C(n16326), .Z(n14151) );
  CMXI2X1 U13223 ( .A0(n18116), .A1(poly1_shifted[177]), .S(n12210), .Z(n14150) );
  COND4CX1 U13224 ( .A(Poly1[155]), .B(Poly1[340]), .C(n14151), .D(n14150), 
        .Z(n9191) );
  CEOXL U13225 ( .A(Poly12[115]), .B(Poly12[26]), .Z(n14154) );
  COND1XL U13226 ( .A(Poly12[122]), .B(n14154), .C(n17613), .Z(n14153) );
  CMXI2X1 U13227 ( .A0(n12013), .A1(poly12_shifted[58]), .S(n12598), .Z(n14152) );
  COND4CX1 U13228 ( .A(n14154), .B(Poly12[122]), .C(n14153), .D(n14152), .Z(
        n10490) );
  COND1XL U13229 ( .A(Poly5[85]), .B(Poly5[120]), .C(n16326), .Z(n14156) );
  CMXI2X1 U13230 ( .A0(n18053), .A1(Poly5[99]), .S(n15403), .Z(n14155) );
  COND4CX1 U13231 ( .A(Poly5[120]), .B(Poly5[85]), .C(n14156), .D(n14155), .Z(
        n11427) );
  COND1XL U13232 ( .A(Poly1[342]), .B(Poly1[157]), .C(n17072), .Z(n14158) );
  CMXI2X1 U13233 ( .A0(n18142), .A1(poly1_shifted[179]), .S(n12210), .Z(n14157) );
  COND4CX1 U13234 ( .A(Poly1[157]), .B(Poly1[342]), .C(n14158), .D(n14157), 
        .Z(n9189) );
  COND1XL U13235 ( .A(Poly0[214]), .B(Poly0[17]), .C(n16702), .Z(n14161) );
  CANR2X1 U13236 ( .A(n18053), .B(n14159), .C(n17500), .D(poly0_shifted[53]), 
        .Z(n14160) );
  COND4CX1 U13237 ( .A(Poly0[17]), .B(Poly0[214]), .C(n14161), .D(n14160), .Z(
        n9542) );
  COND1XL U13238 ( .A(Poly0[212]), .B(Poly0[160]), .C(n17965), .Z(n14163) );
  CANR2X1 U13239 ( .A(n18210), .B(n15960), .C(poly0_shifted[196]), .D(n15671), 
        .Z(n14162) );
  COND4CX1 U13240 ( .A(Poly0[160]), .B(Poly0[212]), .C(n14163), .D(n14162), 
        .Z(n9399) );
  COND1XL U13241 ( .A(Poly13[522]), .B(Poly13[395]), .C(n16702), .Z(n14165) );
  CMXI2X1 U13242 ( .A0(n18249), .A1(poly13_shifted[423]), .S(n17043), .Z(
        n14164) );
  COND4CX1 U13243 ( .A(Poly13[395]), .B(Poly13[522]), .C(n14165), .D(n14164), 
        .Z(n10651) );
  COND1XL U13244 ( .A(Poly6[27]), .B(Poly6[55]), .C(n16919), .Z(n14168) );
  CMXI2X1 U13245 ( .A0(n11986), .A1(Poly6[37]), .S(n14166), .Z(n14167) );
  COND4CX1 U13246 ( .A(Poly6[55]), .B(Poly6[27]), .C(n14168), .D(n14167), .Z(
        n9656) );
  COND1XL U13247 ( .A(Poly13[274]), .B(Poly13[519]), .C(n16326), .Z(n14170) );
  CMXI2X1 U13248 ( .A0(n12010), .A1(poly13_shifted[302]), .S(n17615), .Z(
        n14169) );
  COND4CX1 U13249 ( .A(Poly13[519]), .B(Poly13[274]), .C(n14170), .D(n14169), 
        .Z(n10772) );
  COND1XL U13250 ( .A(Poly1[341]), .B(Poly1[156]), .C(n17466), .Z(n14172) );
  CMXI2X1 U13251 ( .A0(n18138), .A1(poly1_shifted[178]), .S(n12210), .Z(n14171) );
  COND4CX1 U13252 ( .A(Poly1[156]), .B(Poly1[341]), .C(n14172), .D(n14171), 
        .Z(n9190) );
  CANR2X1 U13253 ( .A(n18116), .B(n14505), .C(n17503), .D(Poly0[6]), .Z(n14173) );
  CND2X1 U13254 ( .A(n17642), .B(Poly0[208]), .Z(n14508) );
  CND2X1 U13255 ( .A(n14173), .B(n14508), .Z(n9571) );
  COND1XL U13256 ( .A(Poly0[214]), .B(Poly0[162]), .C(n17965), .Z(n14175) );
  CANR2X1 U13257 ( .A(n18082), .B(n15960), .C(poly0_shifted[198]), .D(n17314), 
        .Z(n14174) );
  COND4CX1 U13258 ( .A(Poly0[162]), .B(Poly0[214]), .C(n14175), .D(n14174), 
        .Z(n9397) );
  COND1XL U13259 ( .A(Poly1[343]), .B(Poly1[205]), .C(n17238), .Z(n14177) );
  CMXI2X1 U13260 ( .A0(n13994), .A1(poly1_shifted[227]), .S(n17053), .Z(n14176) );
  COND4CX1 U13261 ( .A(Poly1[205]), .B(Poly1[343]), .C(n14177), .D(n14176), 
        .Z(n9141) );
  COND1XL U13262 ( .A(Poly0[202]), .B(Poly0[150]), .C(n18047), .Z(n14179) );
  CANR2X1 U13263 ( .A(n18142), .B(n15960), .C(n17314), .D(poly0_shifted[186]), 
        .Z(n14178) );
  COND4CX1 U13264 ( .A(Poly0[150]), .B(Poly0[202]), .C(n14179), .D(n14178), 
        .Z(n9409) );
  CEOXL U13265 ( .A(Poly8[91]), .B(Poly8[12]), .Z(n14182) );
  COND1XL U13266 ( .A(Poly8[93]), .B(n14182), .C(n17285), .Z(n14181) );
  CMXI2X1 U13267 ( .A0(n18095), .A1(poly8_shifted[40]), .S(n12175), .Z(n14180)
         );
  COND4CX1 U13268 ( .A(n14182), .B(Poly8[93]), .C(n14181), .D(n14180), .Z(
        n11375) );
  CEOXL U13269 ( .A(Poly8[85]), .B(Poly8[4]), .Z(n14185) );
  COND1XL U13270 ( .A(Poly8[83]), .B(n14185), .C(n17613), .Z(n14184) );
  CMXI2X1 U13271 ( .A0(n18210), .A1(poly8_shifted[32]), .S(n12175), .Z(n14183)
         );
  COND4CX1 U13272 ( .A(n14185), .B(Poly8[83]), .C(n14184), .D(n14183), .Z(
        n11383) );
  COND1XL U13273 ( .A(Poly8[2]), .B(Poly8[83]), .C(n17398), .Z(n14187) );
  CMXI2X1 U13274 ( .A0(n18167), .A1(Poly8[16]), .S(n12175), .Z(n14186) );
  COND4CX1 U13275 ( .A(Poly8[83]), .B(Poly8[2]), .C(n14187), .D(n14186), .Z(
        n11385) );
  COND1XL U13276 ( .A(Poly3[75]), .B(Poly3[36]), .C(n16372), .Z(n14189) );
  CMXI2X1 U13277 ( .A0(n18210), .A1(Poly3[50]), .S(n17262), .Z(n14188) );
  COND4CX1 U13278 ( .A(Poly3[36]), .B(Poly3[75]), .C(n14189), .D(n14188), .Z(
        n8890) );
  COND1XL U13279 ( .A(Poly0[219]), .B(Poly0[120]), .C(n17705), .Z(n14192) );
  CANR2X1 U13280 ( .A(n12013), .B(n14441), .C(n17671), .D(poly0_shifted[156]), 
        .Z(n14191) );
  COND4CX1 U13281 ( .A(Poly0[120]), .B(Poly0[219]), .C(n14192), .D(n14191), 
        .Z(n9439) );
  COND1XL U13282 ( .A(Poly0[211]), .B(Poly0[112]), .C(n17714), .Z(n14194) );
  CANR2X1 U13283 ( .A(n13428), .B(n14441), .C(n17671), .D(poly0_shifted[148]), 
        .Z(n14193) );
  COND4CX1 U13284 ( .A(Poly0[112]), .B(Poly0[211]), .C(n14194), .D(n14193), 
        .Z(n9447) );
  COND1XL U13285 ( .A(Poly0[114]), .B(Poly0[213]), .C(n17714), .Z(n14196) );
  CANR2X1 U13286 ( .A(n12004), .B(n14441), .C(n17671), .D(poly0_shifted[150]), 
        .Z(n14195) );
  COND4CX1 U13287 ( .A(Poly0[213]), .B(Poly0[114]), .C(n14196), .D(n14195), 
        .Z(n9445) );
  COND1XL U13288 ( .A(Poly0[119]), .B(Poly0[218]), .C(n18234), .Z(n14198) );
  CANR2X1 U13289 ( .A(n18189), .B(n14441), .C(n17671), .D(poly0_shifted[155]), 
        .Z(n14197) );
  COND4CX1 U13290 ( .A(Poly0[218]), .B(Poly0[119]), .C(n14198), .D(n14197), 
        .Z(n9440) );
  COND1XL U13291 ( .A(Poly0[212]), .B(Poly0[113]), .C(n17317), .Z(n14200) );
  CANR2X1 U13292 ( .A(n18053), .B(n14441), .C(n17671), .D(poly0_shifted[149]), 
        .Z(n14199) );
  COND4CX1 U13293 ( .A(Poly0[113]), .B(Poly0[212]), .C(n14200), .D(n14199), 
        .Z(n9446) );
  COND1XL U13294 ( .A(Poly0[210]), .B(Poly0[111]), .C(n17714), .Z(n14202) );
  CANR2X1 U13295 ( .A(n14765), .B(n14441), .C(n17671), .D(poly0_shifted[147]), 
        .Z(n14201) );
  COND4CX1 U13296 ( .A(Poly0[111]), .B(Poly0[210]), .C(n14202), .D(n14201), 
        .Z(n9448) );
  COND1XL U13297 ( .A(Poly0[116]), .B(Poly0[215]), .C(n17508), .Z(n14204) );
  CANR2X1 U13298 ( .A(n14754), .B(n14441), .C(n17671), .D(poly0_shifted[152]), 
        .Z(n14203) );
  COND4CX1 U13299 ( .A(Poly0[215]), .B(Poly0[116]), .C(n14204), .D(n14203), 
        .Z(n9443) );
  COND1XL U13300 ( .A(Poly0[110]), .B(Poly0[209]), .C(n17714), .Z(n14206) );
  CANR2X1 U13301 ( .A(n18108), .B(n14441), .C(n17671), .D(poly0_shifted[146]), 
        .Z(n14205) );
  COND4CX1 U13302 ( .A(Poly0[209]), .B(Poly0[110]), .C(n14206), .D(n14205), 
        .Z(n9449) );
  COND1XL U13303 ( .A(Poly0[214]), .B(Poly0[115]), .C(n17552), .Z(n14208) );
  CANR2X1 U13304 ( .A(n11982), .B(n14441), .C(n17671), .D(poly0_shifted[151]), 
        .Z(n14207) );
  COND4CX1 U13305 ( .A(Poly0[115]), .B(Poly0[214]), .C(n14208), .D(n14207), 
        .Z(n9444) );
  COND1XL U13306 ( .A(Poly3[81]), .B(Poly3[56]), .C(n17527), .Z(n14210) );
  CANR2X1 U13307 ( .A(n14754), .B(n18209), .C(Poly3[70]), .D(n17359), .Z(
        n14209) );
  COND4CX1 U13308 ( .A(Poly3[56]), .B(Poly3[81]), .C(n14210), .D(n14209), .Z(
        n8870) );
  CIVX2 U13309 ( .A(n17259), .Z(n17383) );
  COND1XL U13310 ( .A(Poly3[58]), .B(Poly3[83]), .C(n17383), .Z(n14212) );
  CANR2X1 U13311 ( .A(n18142), .B(n18209), .C(Poly3[72]), .D(n17359), .Z(
        n14211) );
  COND4CX1 U13312 ( .A(Poly3[83]), .B(Poly3[58]), .C(n14212), .D(n14211), .Z(
        n8868) );
  CIVX1 U13313 ( .A(n15168), .Z(n14457) );
  CND2X1 U13314 ( .A(n14213), .B(n11972), .Z(n14979) );
  COND2X1 U13315 ( .A(n14686), .B(n14660), .C(n14979), .D(n15044), .Z(n14215)
         );
  CANR3X1 U13316 ( .A(entrophy[24]), .B(n14457), .C(n14215), .D(n14214), .Z(
        n14237) );
  CND2X1 U13317 ( .A(n13945), .B(datain[6]), .Z(n14685) );
  CND2XL U13318 ( .A(n15206), .B(entrophy[29]), .Z(n14216) );
  CND4X1 U13319 ( .A(n17766), .B(n14685), .C(n14218), .D(n14216), .Z(n14224)
         );
  CNR2X1 U13320 ( .A(n15351), .B(n14886), .Z(n14955) );
  CIVX1 U13321 ( .A(n14955), .Z(n14219) );
  CAN4X1 U13322 ( .A(n14219), .B(n14218), .C(n14217), .D(n15248), .Z(n14220)
         );
  CANR4CX1 U13323 ( .A(n14453), .B(n14451), .C(n14220), .D(n15112), .Z(n14223)
         );
  CND2X1 U13324 ( .A(n17759), .B(datain[3]), .Z(n14987) );
  CND2XL U13325 ( .A(n17495), .B(scrambler[16]), .Z(n14221) );
  COND1XL U13326 ( .A(n15293), .B(n14987), .C(n14221), .Z(n14222) );
  CANR3X1 U13327 ( .A(n15309), .B(n14224), .C(n14223), .D(n14222), .Z(n14236)
         );
  CIVX1 U13328 ( .A(n15006), .Z(n14228) );
  CNR2X1 U13329 ( .A(n14226), .B(n14225), .Z(n14475) );
  CNR2XL U13330 ( .A(n14475), .B(n14866), .Z(n14227) );
  CND2X1 U13331 ( .A(n17759), .B(entrophy[6]), .Z(n15070) );
  CND2X1 U13332 ( .A(n15206), .B(datain[6]), .Z(n14986) );
  CND2X1 U13333 ( .A(n15256), .B(entrophy[25]), .Z(n15140) );
  CND2X1 U13334 ( .A(n11974), .B(datain[0]), .Z(n14704) );
  CND2X1 U13335 ( .A(n15206), .B(entrophy[2]), .Z(n15096) );
  CND2X1 U13336 ( .A(n15256), .B(datain[2]), .Z(n15172) );
  CIVX4 U13337 ( .A(n14230), .Z(n15348) );
  CIVX1 U13338 ( .A(n14231), .Z(n14233) );
  COND3X1 U13339 ( .A(n14237), .B(n14977), .C(n14236), .D(n14235), .Z(n8716)
         );
  CEOXL U13340 ( .A(Poly12[121]), .B(Poly12[62]), .Z(n14240) );
  COND1XL U13341 ( .A(Poly12[122]), .B(n14240), .C(n18234), .Z(n14239) );
  CMXI2X1 U13342 ( .A0(n18160), .A1(poly12_shifted[94]), .S(n12161), .Z(n14238) );
  COND4CX1 U13343 ( .A(n14240), .B(Poly12[122]), .C(n14239), .D(n14238), .Z(
        n10454) );
  CEOXL U13344 ( .A(Poly12[122]), .B(Poly12[63]), .Z(n14243) );
  COND1XL U13345 ( .A(Poly12[123]), .B(n14243), .C(n17538), .Z(n14242) );
  CMXI2X1 U13346 ( .A0(n18206), .A1(poly12_shifted[95]), .S(n12161), .Z(n14241) );
  COND4CX1 U13347 ( .A(n14243), .B(Poly12[123]), .C(n14242), .D(n14241), .Z(
        n10453) );
  COND1XL U13348 ( .A(Poly12[111]), .B(Poly12[51]), .C(n16488), .Z(n14245) );
  CMXI2X1 U13349 ( .A0(n18053), .A1(Poly12[67]), .S(n12161), .Z(n14244) );
  COND4CX1 U13350 ( .A(Poly12[51]), .B(Poly12[111]), .C(n14245), .D(n14244), 
        .Z(n10465) );
  CEOXL U13351 ( .A(Poly12[64]), .B(Poly12[124]), .Z(n14248) );
  COND1XL U13352 ( .A(Poly12[123]), .B(n14248), .C(n18234), .Z(n14247) );
  CMXI2X1 U13353 ( .A0(n18167), .A1(poly12_shifted[96]), .S(n12161), .Z(n14246) );
  COND4CX1 U13354 ( .A(n14248), .B(Poly12[123]), .C(n14247), .D(n14246), .Z(
        n10452) );
  CEOXL U13355 ( .A(Poly12[115]), .B(Poly12[56]), .Z(n14251) );
  COND1XL U13356 ( .A(Poly12[116]), .B(n14251), .C(n17538), .Z(n14250) );
  CMXI2X1 U13357 ( .A0(n18142), .A1(poly12_shifted[88]), .S(n12161), .Z(n14249) );
  COND4CX1 U13358 ( .A(n14251), .B(Poly12[116]), .C(n14250), .D(n14249), .Z(
        n10460) );
  CEOXL U13359 ( .A(Poly12[125]), .B(Poly12[65]), .Z(n14254) );
  COND1XL U13360 ( .A(Poly12[124]), .B(n14254), .C(n17072), .Z(n14253) );
  CMXI2X1 U13361 ( .A0(n13522), .A1(Poly12[81]), .S(n12161), .Z(n14252) );
  COND4CX1 U13362 ( .A(n14254), .B(Poly12[124]), .C(n14253), .D(n14252), .Z(
        n10451) );
  COND1XL U13363 ( .A(Poly1[336]), .B(Poly1[225]), .C(n17156), .Z(n14256) );
  CMXI2X1 U13364 ( .A0(n13028), .A1(poly1_shifted[247]), .S(n12192), .Z(n14255) );
  COND4CX1 U13365 ( .A(Poly1[225]), .B(Poly1[336]), .C(n14256), .D(n14255), 
        .Z(n9121) );
  CIVX2 U13366 ( .A(n17259), .Z(n17334) );
  COND1XL U13367 ( .A(Poly3[73]), .B(Poly3[34]), .C(n17334), .Z(n14258) );
  CMXI2X1 U13368 ( .A0(n18167), .A1(Poly3[48]), .S(n17262), .Z(n14257) );
  COND4CX1 U13369 ( .A(Poly3[34]), .B(Poly3[73]), .C(n14258), .D(n14257), .Z(
        n8892) );
  COND1XL U13370 ( .A(Poly1[342]), .B(Poly1[231]), .C(n17642), .Z(n14260) );
  CMXI2X1 U13371 ( .A0(n18210), .A1(poly1_shifted[253]), .S(n12192), .Z(n14259) );
  COND4CX1 U13372 ( .A(Poly1[231]), .B(Poly1[342]), .C(n14260), .D(n14259), 
        .Z(n9115) );
  COND1XL U13373 ( .A(Poly1[346]), .B(Poly1[235]), .C(n16435), .Z(n14262) );
  CMXI2X1 U13374 ( .A0(n14487), .A1(poly1_shifted[257]), .S(n12192), .Z(n14261) );
  COND4CX1 U13375 ( .A(Poly1[235]), .B(Poly1[346]), .C(n14262), .D(n14261), 
        .Z(n9111) );
  COND1XL U13376 ( .A(Poly1[345]), .B(Poly1[207]), .C(n16583), .Z(n14264) );
  CMXI2X1 U13377 ( .A0(n18095), .A1(poly1_shifted[229]), .S(n17053), .Z(n14263) );
  COND4CX1 U13378 ( .A(Poly1[207]), .B(Poly1[345]), .C(n14264), .D(n14263), 
        .Z(n9139) );
  COND1XL U13379 ( .A(Poly1[337]), .B(Poly1[226]), .C(n17348), .Z(n14266) );
  CMXI2X1 U13380 ( .A0(n18219), .A1(poly1_shifted[248]), .S(n12192), .Z(n14265) );
  COND4CX1 U13381 ( .A(Poly1[226]), .B(Poly1[337]), .C(n14266), .D(n14265), 
        .Z(n9120) );
  COND1XL U13382 ( .A(Poly1[345]), .B(Poly1[234]), .C(n17198), .Z(n14268) );
  CMXI2X1 U13383 ( .A0(n18241), .A1(poly1_shifted[256]), .S(n12192), .Z(n14267) );
  COND4CX1 U13384 ( .A(Poly1[234]), .B(Poly1[345]), .C(n14268), .D(n14267), 
        .Z(n9112) );
  COND1XL U13385 ( .A(Poly1[338]), .B(Poly1[227]), .C(n17198), .Z(n14270) );
  CMXI2X1 U13386 ( .A0(n18160), .A1(poly1_shifted[249]), .S(n12192), .Z(n14269) );
  COND4CX1 U13387 ( .A(Poly1[227]), .B(Poly1[338]), .C(n14270), .D(n14269), 
        .Z(n9119) );
  COND1XL U13388 ( .A(Poly1[340]), .B(Poly1[229]), .C(n17533), .Z(n14272) );
  CMXI2X1 U13389 ( .A0(n18167), .A1(poly1_shifted[251]), .S(n12192), .Z(n14271) );
  COND4CX1 U13390 ( .A(Poly1[229]), .B(Poly1[340]), .C(n14272), .D(n14271), 
        .Z(n9117) );
  COND1XL U13391 ( .A(Poly3[31]), .B(Poly3[70]), .C(n17527), .Z(n14274) );
  CMXI2X1 U13392 ( .A0(n18219), .A1(Poly3[45]), .S(n17262), .Z(n14273) );
  COND4CX1 U13393 ( .A(Poly3[70]), .B(Poly3[31]), .C(n14274), .D(n14273), .Z(
        n8895) );
  CIVX2 U13394 ( .A(n17259), .Z(n16502) );
  COND1XL U13395 ( .A(Poly3[72]), .B(Poly3[33]), .C(n16502), .Z(n14276) );
  CMXI2X1 U13396 ( .A0(n18206), .A1(Poly3[47]), .S(n17262), .Z(n14275) );
  COND4CX1 U13397 ( .A(Poly3[33]), .B(Poly3[72]), .C(n14276), .D(n14275), .Z(
        n8893) );
  COND1XL U13398 ( .A(Poly1[341]), .B(Poly1[230]), .C(n17121), .Z(n14278) );
  CMXI2X1 U13399 ( .A0(n18048), .A1(poly1_shifted[252]), .S(n12192), .Z(n14277) );
  COND4CX1 U13400 ( .A(Poly1[230]), .B(Poly1[341]), .C(n14278), .D(n14277), 
        .Z(n9116) );
  CIVX2 U13401 ( .A(n17259), .Z(n17245) );
  COND1XL U13402 ( .A(Poly2[66]), .B(Poly2[39]), .C(n17245), .Z(n14280) );
  CMXI2X1 U13403 ( .A0(n18176), .A1(Poly2[51]), .S(n17306), .Z(n14279) );
  COND4CX1 U13404 ( .A(Poly2[39]), .B(Poly2[66]), .C(n14280), .D(n14279), .Z(
        n8959) );
  CEOXL U13405 ( .A(Poly3[42]), .B(Poly3[75]), .Z(n14283) );
  CIVX2 U13406 ( .A(n17259), .Z(n17144) );
  COND1XL U13407 ( .A(Poly3[81]), .B(n14283), .C(n17144), .Z(n14282) );
  CMXI2X1 U13408 ( .A0(n13994), .A1(Poly3[56]), .S(n17262), .Z(n14281) );
  COND4CX1 U13409 ( .A(n14283), .B(Poly3[81]), .C(n14282), .D(n14281), .Z(
        n8884) );
  CEOX1 U13410 ( .A(Poly12[121]), .B(Poly12[61]), .Z(n14288) );
  CND2X1 U13411 ( .A(n14284), .B(n14288), .Z(n14286) );
  CMXI2X1 U13412 ( .A0(n18219), .A1(poly12_shifted[93]), .S(n12161), .Z(n14285) );
  COND3X1 U13413 ( .A(n14288), .B(n14287), .C(n14286), .D(n14285), .Z(n10455)
         );
  CEOX1 U13414 ( .A(Poly12[54]), .B(Poly12[114]), .Z(n14291) );
  CND2X1 U13415 ( .A(n14292), .B(n14291), .Z(n14290) );
  CMXI2X1 U13416 ( .A0(n14754), .A1(poly12_shifted[86]), .S(n12161), .Z(n14289) );
  COND3X1 U13417 ( .A(n14291), .B(n14295), .C(n14290), .D(n14289), .Z(n10462)
         );
  CEOX1 U13418 ( .A(Poly12[112]), .B(Poly12[53]), .Z(n14296) );
  CND2X1 U13419 ( .A(n14292), .B(n14296), .Z(n14294) );
  CMXI2X1 U13420 ( .A0(n11992), .A1(poly12_shifted[85]), .S(n12161), .Z(n14293) );
  COND3X1 U13421 ( .A(n14296), .B(n14295), .C(n14294), .D(n14293), .Z(n10463)
         );
  COND1XL U13422 ( .A(Poly3[74]), .B(Poly3[35]), .C(n16540), .Z(n14299) );
  CMXI2X1 U13423 ( .A0(n14297), .A1(Poly3[49]), .S(n17262), .Z(n14298) );
  COND4CX1 U13424 ( .A(Poly3[35]), .B(Poly3[74]), .C(n14299), .D(n14298), .Z(
        n8891) );
  CND2X1 U13425 ( .A(n14300), .B(Poly11[24]), .Z(n14302) );
  CMXI2X1 U13426 ( .A0(n18138), .A1(Poly11[39]), .S(n17683), .Z(n14301) );
  COND3X1 U13427 ( .A(Poly11[24]), .B(n14303), .C(n14302), .D(n14301), .Z(
        n11150) );
  COND1XL U13428 ( .A(Poly14[292]), .B(Poly14[172]), .C(n17290), .Z(n14305) );
  COND4CX1 U13429 ( .A(Poly14[172]), .B(Poly14[292]), .C(n14305), .D(n14304), 
        .Z(n10217) );
  COND1XL U13430 ( .A(Poly14[290]), .B(Poly14[170]), .C(n17535), .Z(n14307) );
  CMXI2X1 U13431 ( .A0(n18095), .A1(poly14_shifted[202]), .S(n13129), .Z(
        n14306) );
  COND4CX1 U13432 ( .A(Poly14[170]), .B(Poly14[290]), .C(n14307), .D(n14306), 
        .Z(n10219) );
  COND1XL U13433 ( .A(Poly14[289]), .B(Poly14[169]), .C(n17755), .Z(n14309) );
  CMXI2X1 U13434 ( .A0(n18249), .A1(poly14_shifted[201]), .S(n13129), .Z(
        n14308) );
  COND4CX1 U13435 ( .A(Poly14[169]), .B(Poly14[289]), .C(n14309), .D(n14308), 
        .Z(n10220) );
  COND1XL U13436 ( .A(Poly6[46]), .B(Poly6[10]), .C(n17401), .Z(n14312) );
  CMXI2X1 U13437 ( .A0(n18082), .A1(Poly6[20]), .S(n14310), .Z(n14311) );
  COND4CX1 U13438 ( .A(Poly6[10]), .B(Poly6[46]), .C(n14312), .D(n14311), .Z(
        n9673) );
  COND1XL U13439 ( .A(Poly1[344]), .B(Poly1[233]), .C(n16312), .Z(n14314) );
  CMXI2X1 U13440 ( .A0(n18082), .A1(poly1_shifted[255]), .S(n12192), .Z(n14313) );
  COND4CX1 U13441 ( .A(Poly1[233]), .B(Poly1[344]), .C(n14314), .D(n14313), 
        .Z(n9113) );
  COND1XL U13442 ( .A(n14317), .B(dataselector[19]), .C(n16919), .Z(n14316) );
  CANR2X1 U13443 ( .A(n18095), .B(n17832), .C(dataselector[26]), .D(n16410), 
        .Z(n14315) );
  COND4CX1 U13444 ( .A(dataselector[19]), .B(n14317), .C(n14316), .D(n14315), 
        .Z(n8769) );
  CND2X1 U13445 ( .A(n15361), .B(poly5_shifted[55]), .Z(n14319) );
  CND2X1 U13446 ( .A(n16644), .B(poly5_shifted[41]), .Z(n14318) );
  COND3X1 U13447 ( .A(n17935), .B(n17208), .C(n14319), .D(n14318), .Z(n11485)
         );
  CNR2X1 U13448 ( .A(Poly15[16]), .B(n18050), .Z(n14320) );
  CENX1 U13449 ( .A(n14321), .B(n14320), .Z(n14322) );
  COND1XL U13450 ( .A(Poly9[106]), .B(Poly9[14]), .C(n17401), .Z(n14325) );
  CMXI2X1 U13451 ( .A0(n18249), .A1(Poly9[25]), .S(n17731), .Z(n14324) );
  COND4CX1 U13452 ( .A(Poly9[14]), .B(Poly9[106]), .C(n14325), .D(n14324), .Z(
        n11280) );
  CEOXL U13453 ( .A(Poly9[109]), .B(Poly9[20]), .Z(n14328) );
  COND1XL U13454 ( .A(Poly9[112]), .B(n14328), .C(n17634), .Z(n14327) );
  CMXI2X1 U13455 ( .A0(n14436), .A1(poly9_shifted[42]), .S(n17731), .Z(n14326)
         );
  COND4CX1 U13456 ( .A(n14328), .B(Poly9[112]), .C(n14327), .D(n14326), .Z(
        n11274) );
  COND1XL U13457 ( .A(Poly3[77]), .B(Poly3[52]), .C(n17343), .Z(n14330) );
  CANR2X1 U13458 ( .A(n13428), .B(n18209), .C(n17359), .D(poly3_shifted[80]), 
        .Z(n14329) );
  COND4CX1 U13459 ( .A(Poly3[52]), .B(Poly3[77]), .C(n14330), .D(n14329), .Z(
        n8874) );
  COND1XL U13460 ( .A(Poly3[80]), .B(Poly3[55]), .C(n17099), .Z(n14332) );
  CANR2X1 U13461 ( .A(n11996), .B(n18209), .C(n17359), .D(poly3_shifted[83]), 
        .Z(n14331) );
  COND4CX1 U13462 ( .A(Poly3[55]), .B(Poly3[80]), .C(n14332), .D(n14331), .Z(
        n8871) );
  COND1XL U13463 ( .A(Poly3[76]), .B(Poly3[51]), .C(n17121), .Z(n14334) );
  CANR2X1 U13464 ( .A(n14361), .B(n18209), .C(n17359), .D(poly3_shifted[79]), 
        .Z(n14333) );
  COND4CX1 U13465 ( .A(Poly3[51]), .B(Poly3[76]), .C(n14334), .D(n14333), .Z(
        n8875) );
  COND1XL U13466 ( .A(Poly3[53]), .B(Poly3[78]), .C(n17466), .Z(n14336) );
  CANR2X1 U13467 ( .A(n18053), .B(n18209), .C(n17359), .D(poly3_shifted[81]), 
        .Z(n14335) );
  COND4CX1 U13468 ( .A(Poly3[78]), .B(Poly3[53]), .C(n14336), .D(n14335), .Z(
        n8873) );
  CND2XL U13469 ( .A(poly0_shifted[192]), .B(n15671), .Z(n14339) );
  CAN2X1 U13470 ( .A(n17538), .B(n14337), .Z(n14504) );
  COND4CX1 U13471 ( .A(n14504), .B(Poly0[156]), .C(n18160), .D(n15672), .Z(
        n14338) );
  COND3X1 U13472 ( .A(Poly0[156]), .B(n14508), .C(n14339), .D(n14338), .Z(
        n9403) );
  CIVX2 U13473 ( .A(n15880), .Z(n16276) );
  COND4CXL U13474 ( .A(Poly0[109]), .B(n14504), .C(n12003), .D(n16276), .Z(
        n14341) );
  CND2X1 U13475 ( .A(n15880), .B(poly0_shifted[145]), .Z(n14340) );
  COND3X1 U13476 ( .A(Poly0[109]), .B(n14508), .C(n14341), .D(n14340), .Z(
        n9450) );
  COND1XL U13477 ( .A(Poly7[402]), .B(Poly7[236]), .C(n17538), .Z(n14343) );
  CMXI2X1 U13478 ( .A0(n13994), .A1(poly7_shifted[260]), .S(n17574), .Z(n14342) );
  COND4CX1 U13479 ( .A(Poly7[236]), .B(Poly7[402]), .C(n14343), .D(n14342), 
        .Z(n9856) );
  COND1XL U13480 ( .A(Poly7[406]), .B(Poly7[240]), .C(n17290), .Z(n14345) );
  COND4CX1 U13481 ( .A(Poly7[240]), .B(Poly7[406]), .C(n14345), .D(n14344), 
        .Z(n9852) );
  COND1XL U13482 ( .A(\dataselector_shifted[0] ), .B(Poly7[238]), .C(n18234), 
        .Z(n14347) );
  CMXI2X1 U13483 ( .A0(n18095), .A1(poly7_shifted[262]), .S(n17574), .Z(n14346) );
  COND4CX1 U13484 ( .A(Poly7[238]), .B(\dataselector_shifted[0] ), .C(n14347), 
        .D(n14346), .Z(n9854) );
  CENX1 U13485 ( .A(Poly15[24]), .B(Poly15[50]), .Z(n14348) );
  CENX1 U13486 ( .A(Poly15[56]), .B(n14348), .Z(n14351) );
  COND1XL U13487 ( .A(Poly15[57]), .B(n14351), .C(n17094), .Z(n14350) );
  CMXI2X1 U13488 ( .A0(n18138), .A1(poly15_shifted[54]), .S(n17376), .Z(n14349) );
  COND4CX1 U13489 ( .A(n14351), .B(Poly15[57]), .C(n14350), .D(n14349), .Z(
        n9598) );
  COND1XL U13490 ( .A(Poly15[55]), .B(Poly15[29]), .C(n17504), .Z(n14353) );
  CMXI2X1 U13491 ( .A0(n13028), .A1(poly15_shifted[59]), .S(n17376), .Z(n14352) );
  COND4CX1 U13492 ( .A(Poly15[29]), .B(Poly15[55]), .C(n14353), .D(n14352), 
        .Z(n9593) );
  CIVX1 U13493 ( .A(Poly5[119]), .Z(n15413) );
  CIVX1 U13494 ( .A(Poly5[84]), .Z(n16006) );
  CND2X1 U13495 ( .A(n15413), .B(n16006), .Z(n14357) );
  CND2X1 U13496 ( .A(n17203), .B(n14357), .Z(n14359) );
  CMXI2X1 U13497 ( .A0(n12415), .A1(Poly5[98]), .S(n15403), .Z(n14358) );
  COND4CX1 U13498 ( .A(Poly5[84]), .B(Poly5[119]), .C(n14359), .D(n14358), .Z(
        n11428) );
  CIVXL U13499 ( .A(Poly13[520]), .Z(n14360) );
  CIVXL U13500 ( .A(Poly13[515]), .Z(n14362) );
  CIVXL U13501 ( .A(Poly13[521]), .Z(n14363) );
  CIVXL U13502 ( .A(Poly1[345]), .Z(n14364) );
  COND1XL U13503 ( .A(Poly13[517]), .B(Poly13[158]), .C(n17504), .Z(n14366) );
  CMXI2X1 U13504 ( .A0(n13028), .A1(poly13_shifted[186]), .S(n13014), .Z(
        n14365) );
  COND4CX1 U13505 ( .A(Poly13[158]), .B(Poly13[517]), .C(n14366), .D(n14365), 
        .Z(n10888) );
  COND1XL U13506 ( .A(Poly1[343]), .B(Poly1[60]), .C(n17266), .Z(n14368) );
  CMXI2X1 U13507 ( .A0(n18138), .A1(poly1_shifted[82]), .S(n12012), .Z(n14367)
         );
  COND4CX1 U13508 ( .A(Poly1[60]), .B(Poly1[343]), .C(n14368), .D(n14367), .Z(
        n9286) );
  CND2XL U13509 ( .A(n17959), .B(scrambler[29]), .Z(n14373) );
  CIVX1 U13510 ( .A(n14373), .Z(n14380) );
  CND3XL U13511 ( .A(n14369), .B(n14672), .C(entrophy[8]), .Z(n14371) );
  CNR2X1 U13512 ( .A(n14969), .B(n14926), .Z(n15020) );
  CIVX2 U13513 ( .A(n15020), .Z(n14410) );
  CND2X1 U13514 ( .A(n15319), .B(entrophy[4]), .Z(n15136) );
  CND2X1 U13515 ( .A(n14540), .B(entrophy[30]), .Z(n14901) );
  CND8X1 U13516 ( .A(n14371), .B(n14866), .C(n14370), .D(n14410), .E(n15024), 
        .F(n15136), .G(n14901), .H(n15060), .Z(n14379) );
  CNR2X1 U13517 ( .A(n12018), .B(n17808), .Z(n15296) );
  CAN2X1 U13518 ( .A(n15206), .B(entrophy[9]), .Z(n15058) );
  CNR4X1 U13519 ( .A(n15296), .B(n15058), .C(n15099), .D(n14372), .Z(n14377)
         );
  CAN4X1 U13520 ( .A(n14558), .B(n14652), .C(n14374), .D(n14373), .Z(n14376)
         );
  CND4X1 U13521 ( .A(n14377), .B(n14376), .C(n14375), .D(n15136), .Z(n14378)
         );
  COND3X1 U13522 ( .A(n17804), .B(n14380), .C(n14379), .D(n14378), .Z(n14391)
         );
  CANR2X1 U13523 ( .A(n17770), .B(entrophy[11]), .C(datain[0]), .D(n14976), 
        .Z(n14381) );
  CANR4CX1 U13524 ( .A(n15229), .B(n15332), .C(n14381), .D(n12535), .Z(n14382)
         );
  CND2X1 U13525 ( .A(n12019), .B(entrophy[3]), .Z(n15217) );
  COND3X1 U13526 ( .A(n15300), .B(n14226), .C(n14383), .D(n15217), .Z(n14386)
         );
  CNR2X1 U13527 ( .A(n15283), .B(n14453), .Z(n15311) );
  COND3X1 U13528 ( .A(n14387), .B(n12520), .C(n14892), .D(n14384), .Z(n14385)
         );
  CNR2X1 U13529 ( .A(n14981), .B(n14387), .Z(n15072) );
  CND3XL U13530 ( .A(n14558), .B(n15172), .C(n14388), .Z(n14389) );
  CND2XL U13531 ( .A(n14392), .B(entrophy[15]), .Z(n15148) );
  COND1XL U13532 ( .A(n15339), .B(n14393), .C(n15148), .Z(n15109) );
  CIVXL U13533 ( .A(n15109), .Z(n14394) );
  COND3X1 U13534 ( .A(n14394), .B(n14538), .C(n15190), .D(n14417), .Z(n14407)
         );
  CAN2X1 U13535 ( .A(n14826), .B(entrophy[7]), .Z(n15318) );
  CNR2X1 U13536 ( .A(n14395), .B(n14687), .Z(n15111) );
  CIVX1 U13537 ( .A(n15111), .Z(n15076) );
  CNR3X1 U13538 ( .A(n15076), .B(n14396), .C(n15001), .Z(n14548) );
  COND1XL U13539 ( .A(n15318), .B(n14548), .C(n15309), .Z(n14404) );
  CNR2X1 U13540 ( .A(n14397), .B(n15293), .Z(n14402) );
  CNR2X1 U13541 ( .A(n12055), .B(n17784), .Z(n14398) );
  CND2X1 U13542 ( .A(n14857), .B(n14398), .Z(n14400) );
  CND2XL U13543 ( .A(n17826), .B(scrambler[0]), .Z(n14399) );
  CND2X1 U13544 ( .A(n14400), .B(n14399), .Z(n14401) );
  CNR2X1 U13545 ( .A(n14402), .B(n14401), .Z(n14403) );
  CND2X1 U13546 ( .A(n14404), .B(n14403), .Z(n14406) );
  CIVX2 U13547 ( .A(n14877), .Z(n17800) );
  CANR4CX1 U13548 ( .A(n14226), .B(n17800), .C(n14958), .D(n14659), .Z(n14405)
         );
  CANR3X1 U13549 ( .A(n15145), .B(n14407), .C(n14406), .D(n14405), .Z(n14429)
         );
  CIVX1 U13550 ( .A(n14568), .Z(n14408) );
  CND3XL U13551 ( .A(n14408), .B(entrophy[23]), .C(n15798), .Z(n15008) );
  CNR2X1 U13552 ( .A(n14409), .B(n15021), .Z(n14411) );
  CND4X1 U13553 ( .A(n15008), .B(n14411), .C(n17766), .D(n14410), .Z(n14412)
         );
  CANR2X1 U13554 ( .A(n14413), .B(n17804), .C(n15314), .D(n14412), .Z(n14428)
         );
  CND2X1 U13555 ( .A(n14826), .B(datain[5]), .Z(n15061) );
  CND2X1 U13556 ( .A(n15061), .B(n14414), .Z(n15003) );
  CND4X1 U13557 ( .A(n14690), .B(n14417), .C(n14416), .D(n14415), .Z(n14419)
         );
  CND2X1 U13558 ( .A(n17776), .B(entrophy[27]), .Z(n14893) );
  COND11X1 U13559 ( .A(n15003), .B(n14419), .C(n14418), .D(n12216), .Z(n14427)
         );
  COND4CX1 U13560 ( .A(n15075), .B(n14935), .C(n14545), .D(n14420), .Z(n14425)
         );
  CIVXL U13561 ( .A(n14880), .Z(n14423) );
  CANR2XL U13562 ( .A(n15274), .B(entrophy[25]), .C(n14879), .D(n15043), .Z(
        n14422) );
  COND3X1 U13563 ( .A(n14644), .B(n14423), .C(n14422), .D(n14421), .Z(n14424)
         );
  COND1X1 U13564 ( .A(n14425), .B(n14424), .C(n14868), .Z(n14426) );
  CND4X1 U13565 ( .A(n14429), .B(n14428), .C(n14427), .D(n14426), .Z(n8700) );
  COND1XL U13566 ( .A(Poly4[58]), .B(n15651), .C(n17206), .Z(n14431) );
  CMXI2X1 U13567 ( .A0(n13028), .A1(poly4_shifted[29]), .S(n18230), .Z(n14430)
         );
  COND4CX1 U13568 ( .A(n15651), .B(Poly4[58]), .C(n14431), .D(n14430), .Z(
        n8844) );
  COND1XL U13569 ( .A(Poly4[58]), .B(Poly4[60]), .C(n17203), .Z(n14433) );
  CMXI2X1 U13570 ( .A0(n18160), .A1(poly4_shifted[31]), .S(n18230), .Z(n14432)
         );
  COND4CX1 U13571 ( .A(Poly4[60]), .B(Poly4[58]), .C(n14433), .D(n14432), .Z(
        n8842) );
  COND1XL U13572 ( .A(Poly7[403]), .B(Poly7[23]), .C(n16702), .Z(n14435) );
  CMXI2X1 U13573 ( .A0(n18053), .A1(poly7_shifted[47]), .S(n12170), .Z(n14434)
         );
  COND4CX1 U13574 ( .A(Poly7[23]), .B(Poly7[403]), .C(n14435), .D(n14434), .Z(
        n10069) );
  CIVX2 U13575 ( .A(n15673), .Z(n17352) );
  COND1XL U13576 ( .A(Poly14[295]), .B(Poly14[175]), .C(n17352), .Z(n14438) );
  CMXI2X1 U13577 ( .A0(n14436), .A1(poly14_shifted[207]), .S(n13129), .Z(
        n14437) );
  COND4CX1 U13578 ( .A(Poly14[175]), .B(Poly14[295]), .C(n14438), .D(n14437), 
        .Z(n10214) );
  CND2XL U13579 ( .A(n17755), .B(poly9_shifted[52]), .Z(n14440) );
  CND2X1 U13580 ( .A(n13351), .B(poly9_shifted[63]), .Z(n14439) );
  COND4CX1 U13581 ( .A(n14440), .B(n17707), .C(n13351), .D(n14439), .Z(n11253)
         );
  COND1XL U13582 ( .A(Poly0[217]), .B(Poly0[118]), .C(n16502), .Z(n14443) );
  CANR2X1 U13583 ( .A(n18142), .B(n14441), .C(n17671), .D(poly0_shifted[154]), 
        .Z(n14442) );
  COND4CX1 U13584 ( .A(Poly0[118]), .B(Poly0[217]), .C(n14443), .D(n14442), 
        .Z(n9441) );
  COND1XL U13585 ( .A(Poly7[400]), .B(Poly7[20]), .C(n17998), .Z(n14445) );
  CMXI2X1 U13586 ( .A0(n12010), .A1(poly7_shifted[44]), .S(n12170), .Z(n14444)
         );
  COND4CX1 U13587 ( .A(Poly7[20]), .B(Poly7[400]), .C(n14445), .D(n14444), .Z(
        n10072) );
  COND1XL U13588 ( .A(n14448), .B(dataselector[41]), .C(n18047), .Z(n14447) );
  CANR2X1 U13589 ( .A(n18167), .B(n18248), .C(n15710), .D(dataselector[48]), 
        .Z(n14446) );
  COND4CX1 U13590 ( .A(dataselector[41]), .B(n14448), .C(n14447), .D(n14446), 
        .Z(n8747) );
  COND1XL U13591 ( .A(Poly5[115]), .B(Poly5[93]), .C(n17449), .Z(n14450) );
  CMXI2X1 U13592 ( .A0(n16381), .A1(poly5_shifted[121]), .S(n15403), .Z(n14449) );
  COND4CX1 U13593 ( .A(Poly5[93]), .B(Poly5[115]), .C(n14450), .D(n14449), .Z(
        n11419) );
  CIVX2 U13594 ( .A(n14451), .Z(n15074) );
  CANR1XL U13595 ( .A(n14866), .B(n15074), .C(n14976), .Z(n14452) );
  CNR3X1 U13596 ( .A(n12520), .B(n14453), .C(n17800), .Z(n14456) );
  CND2X1 U13597 ( .A(n14454), .B(entrophy[17]), .Z(n17765) );
  COND2X1 U13598 ( .A(n14808), .B(n15075), .C(dataselector[14]), .D(n17765), 
        .Z(n14455) );
  CANR3X1 U13599 ( .A(n14457), .B(datain[5]), .C(n14456), .D(n14455), .Z(
        n14464) );
  CNR2X1 U13600 ( .A(n17759), .B(entrophy[26]), .Z(n14458) );
  CANR3X1 U13601 ( .A(n14967), .B(n14850), .C(n14458), .D(n14652), .Z(n14461)
         );
  CND2X1 U13602 ( .A(n14695), .B(entrophy[31]), .Z(n14779) );
  CND2XL U13603 ( .A(n17829), .B(scrambler[14]), .Z(n14462) );
  CND3XL U13604 ( .A(n17767), .B(n14633), .C(datain[3]), .Z(n14459) );
  COND3X1 U13605 ( .A(n14779), .B(n17785), .C(n14462), .D(n14459), .Z(n14460)
         );
  CANR1XL U13606 ( .A(n14970), .B(n14461), .C(n14460), .Z(n14463) );
  CANR2X1 U13607 ( .A(n14464), .B(n14463), .C(n12535), .D(n14462), .Z(n14480)
         );
  CND2X1 U13608 ( .A(n17770), .B(entrophy[12]), .Z(n15041) );
  CNR2X1 U13609 ( .A(n12535), .B(n14871), .Z(n14661) );
  CNR2X1 U13610 ( .A(n14977), .B(n14465), .Z(n14466) );
  CNR2IX1 U13611 ( .B(n14466), .A(n15335), .Z(n14467) );
  CANR1XL U13612 ( .A(n15043), .B(n14661), .C(n14467), .Z(n14468) );
  COND1XL U13613 ( .A(n14645), .B(n15041), .C(n14468), .Z(n14479) );
  CND2X1 U13614 ( .A(n11974), .B(entrophy[20]), .Z(n14583) );
  CAN4X1 U13615 ( .A(n14470), .B(n14583), .C(n15345), .D(n14469), .Z(n14477)
         );
  CNR2X1 U13616 ( .A(n14969), .B(n14471), .Z(n15255) );
  CNR2X1 U13617 ( .A(n12459), .B(n14659), .Z(n17769) );
  CNR2X1 U13618 ( .A(n14473), .B(n14795), .Z(n15023) );
  CNR8X1 U13619 ( .A(n14475), .B(n15021), .C(n15255), .D(n14823), .E(n15058), 
        .F(n17769), .G(n14474), .H(n15023), .Z(n14476) );
  COND2X1 U13620 ( .A(n14477), .B(n12055), .C(n14476), .D(n17778), .Z(n14478)
         );
  COR4X1 U13621 ( .A(n14481), .B(n14480), .C(n14479), .D(n14478), .Z(n8714) );
  COND1XL U13622 ( .A(Poly4[41]), .B(n14484), .C(n16540), .Z(n14483) );
  CMXI2X1 U13623 ( .A0(n18095), .A1(Poly4[58]), .S(n12153), .Z(n14482) );
  COND4CX1 U13624 ( .A(n14484), .B(Poly4[41]), .C(n14483), .D(n14482), .Z(
        n8798) );
  CEOX1 U13625 ( .A(Poly4[56]), .B(n14485), .Z(n14486) );
  CENX1 U13626 ( .A(n15640), .B(n14486), .Z(n14490) );
  CIVX2 U13627 ( .A(n15673), .Z(n16540) );
  COND1XL U13628 ( .A(Poly4[37]), .B(n14490), .C(n16540), .Z(n14489) );
  CMXI2X1 U13629 ( .A0(n14487), .A1(Poly4[54]), .S(n12153), .Z(n14488) );
  COND4CX1 U13630 ( .A(n14490), .B(Poly4[37]), .C(n14489), .D(n14488), .Z(
        n8802) );
  CIVX2 U13631 ( .A(n15673), .Z(n17523) );
  COND1XL U13632 ( .A(Poly4[39]), .B(n14493), .C(n17523), .Z(n14492) );
  CMXI2X1 U13633 ( .A0(n13994), .A1(Poly4[56]), .S(n12153), .Z(n14491) );
  COND4CX1 U13634 ( .A(n14493), .B(Poly4[39]), .C(n14492), .D(n14491), .Z(
        n8800) );
  COND1XL U13635 ( .A(Poly0[210]), .B(Poly0[13]), .C(n17965), .Z(n14495) );
  CANR2X1 U13636 ( .A(n14436), .B(n14505), .C(n17503), .D(poly0_shifted[49]), 
        .Z(n14494) );
  COND4CX1 U13637 ( .A(Poly0[13]), .B(Poly0[210]), .C(n14495), .D(n14494), .Z(
        n9546) );
  COND1XL U13638 ( .A(Poly0[202]), .B(Poly0[5]), .C(n17178), .Z(n14497) );
  CANR2X1 U13639 ( .A(n11999), .B(n14505), .C(n17503), .D(poly0_shifted[41]), 
        .Z(n14496) );
  COND4CX1 U13640 ( .A(Poly0[5]), .B(Poly0[202]), .C(n14497), .D(n14496), .Z(
        n9554) );
  COND1XL U13641 ( .A(Poly0[207]), .B(Poly0[10]), .C(n16427), .Z(n14499) );
  CANR2X1 U13642 ( .A(n12007), .B(n14505), .C(n17503), .D(poly0_shifted[46]), 
        .Z(n14498) );
  COND4CX1 U13643 ( .A(Poly0[10]), .B(Poly0[207]), .C(n14499), .D(n14498), .Z(
        n9549) );
  COND1XL U13644 ( .A(Poly0[203]), .B(Poly0[6]), .C(n16326), .Z(n14501) );
  CANR2X1 U13645 ( .A(n13994), .B(n14505), .C(n17503), .D(poly0_shifted[42]), 
        .Z(n14500) );
  COND4CX1 U13646 ( .A(Poly0[6]), .B(Poly0[203]), .C(n14501), .D(n14500), .Z(
        n9553) );
  COND1XL U13647 ( .A(Poly0[204]), .B(Poly0[7]), .C(n17705), .Z(n14503) );
  CANR2X1 U13648 ( .A(n18249), .B(n14505), .C(n17503), .D(poly0_shifted[43]), 
        .Z(n14502) );
  COND4CX1 U13649 ( .A(Poly0[7]), .B(Poly0[204]), .C(n14503), .D(n14502), .Z(
        n9552) );
  CND2X1 U13650 ( .A(n14504), .B(Poly0[11]), .Z(n14507) );
  CANR2X1 U13651 ( .A(n18228), .B(n14505), .C(n17503), .D(poly0_shifted[47]), 
        .Z(n14506) );
  COND3X1 U13652 ( .A(Poly0[11]), .B(n14508), .C(n14507), .D(n14506), .Z(n9548) );
  COND1XL U13653 ( .A(Poly7[403]), .B(Poly7[237]), .C(n17266), .Z(n14510) );
  CMXI2X1 U13654 ( .A0(n18249), .A1(poly7_shifted[261]), .S(n17574), .Z(n14509) );
  COND4CX1 U13655 ( .A(Poly7[237]), .B(Poly7[403]), .C(n14510), .D(n14509), 
        .Z(n9855) );
  CND2XL U13656 ( .A(n17755), .B(poly9_shifted[53]), .Z(n14512) );
  CND2X1 U13657 ( .A(n13351), .B(poly9_shifted[64]), .Z(n14511) );
  COND4CX1 U13658 ( .A(n14512), .B(n17036), .C(n13351), .D(n14511), .Z(n11252)
         );
  CND2X1 U13659 ( .A(n18044), .B(poly15_shifted[16]), .Z(n14513) );
  COND4CX1 U13660 ( .A(n18040), .B(n17697), .C(n18044), .D(n14513), .Z(n9636)
         );
  CND2X1 U13661 ( .A(n18044), .B(Poly15[13]), .Z(n14514) );
  COND4CX1 U13662 ( .A(n17065), .B(n14515), .C(n18044), .D(n14514), .Z(n9624)
         );
  CANR2XL U13663 ( .A(Poly2[68]), .B(n16863), .C(n16860), .D(poly9_shifted[14]), .Z(n14520) );
  CANR2X1 U13664 ( .A(n16843), .B(poly6_shifted[17]), .C(n14516), .D(n16840), 
        .Z(n14519) );
  CANR2X1 U13665 ( .A(n16850), .B(poly7_shifted[322]), .C(n16852), .D(
        poly6_shifted[18]), .Z(n14518) );
  CANR2X1 U13666 ( .A(n12067), .B(Poly4[48]), .C(n16874), .D(poly3_shifted[15]), .Z(n14517) );
  CAN4X1 U13667 ( .A(n14520), .B(n14519), .C(n14518), .D(n14517), .Z(n14536)
         );
  CANR2X1 U13668 ( .A(n16864), .B(poly9_shifted[49]), .C(n16872), .D(
        poly5_shifted[33]), .Z(n14524) );
  CANR2X1 U13669 ( .A(n16855), .B(Poly6[17]), .C(Poly4[21]), .D(n16849), .Z(
        n14523) );
  CANR2X1 U13670 ( .A(n16867), .B(poly10_shifted[19]), .C(n16851), .D(
        poly14_shifted[264]), .Z(n14522) );
  CANR2X1 U13671 ( .A(n12071), .B(Poly11[36]), .C(n16841), .D(
        poly9_shifted[108]), .Z(n14521) );
  CAN4X1 U13672 ( .A(n14524), .B(n14523), .C(n14522), .D(n14521), .Z(n14535)
         );
  CANR2X1 U13673 ( .A(n16844), .B(Poly6[51]), .C(n16838), .D(n17938), .Z(
        n14528) );
  CIVXL U13674 ( .A(n14525), .Z(n14526) );
  CANR2X1 U13675 ( .A(Poly3[77]), .B(n16865), .C(n14526), .D(n16861), .Z(
        n14527) );
  CANR2X1 U13676 ( .A(n16875), .B(Poly15[17]), .C(n16866), .D(Poly10[11]), .Z(
        n14532) );
  CANR2X1 U13677 ( .A(n16842), .B(Poly15[24]), .C(n16854), .D(Poly14[210]), 
        .Z(n14531) );
  CANR2X1 U13678 ( .A(n16876), .B(poly4_shifted[19]), .C(n16862), .D(
        poly7_shifted[158]), .Z(n14530) );
  CANR2X1 U13679 ( .A(n16873), .B(Poly2[26]), .C(n16853), .D(poly9_shifted[22]), .Z(n14529) );
  CAN4X1 U13680 ( .A(n14532), .B(n14531), .C(n14530), .D(n14529), .Z(n14533)
         );
  CND4X1 U13681 ( .A(n14536), .B(n14535), .C(n14534), .D(n14533), .Z(n14537)
         );
  CAOR2X2 U13682 ( .A(polydata[9]), .B(n15673), .C(n14537), .D(n16886), .Z(
        n8693) );
  CANR1X1 U13683 ( .A(scrambler[1]), .B(n17744), .C(n14539), .Z(n14543) );
  CND3XL U13684 ( .A(n15034), .B(n14868), .C(entrophy[10]), .Z(n14542) );
  CND2X1 U13685 ( .A(n14540), .B(datain[1]), .Z(n14656) );
  COR2X1 U13686 ( .A(n14656), .B(n17763), .Z(n14541) );
  CND3X1 U13687 ( .A(n14543), .B(n14542), .C(n14541), .Z(n14544) );
  CNR2X1 U13688 ( .A(n15283), .B(n14545), .Z(n14587) );
  CNR2X1 U13689 ( .A(n14546), .B(n14561), .Z(n15131) );
  COR4X1 U13690 ( .A(n14587), .B(n14548), .C(n15131), .D(n14547), .Z(n14556)
         );
  CND2X1 U13691 ( .A(n17792), .B(entrophy[22]), .Z(n14960) );
  CNR2X1 U13692 ( .A(n14969), .B(n14567), .Z(n15213) );
  CANR2X1 U13693 ( .A(n15312), .B(n14868), .C(n15346), .D(n15213), .Z(n14551)
         );
  CND2XL U13694 ( .A(n17774), .B(entrophy[15]), .Z(n14550) );
  COR2XL U13695 ( .A(n14888), .B(n15112), .Z(n14549) );
  CND3XL U13696 ( .A(n14551), .B(n14550), .C(n14549), .Z(n14555) );
  CND2X1 U13697 ( .A(n15319), .B(entrophy[18]), .Z(n14552) );
  CND3XL U13698 ( .A(n15035), .B(dataselector[21]), .C(entrophy[14]), .Z(
        n14859) );
  CND2X1 U13699 ( .A(n14552), .B(n14859), .Z(n14571) );
  CIVXL U13700 ( .A(n14571), .Z(n14553) );
  CANR11X1 U13701 ( .A(n14553), .B(n14925), .C(n15009), .D(n17800), .Z(n14554)
         );
  CANR3X1 U13702 ( .A(n12216), .B(n14556), .C(n14555), .D(n14554), .Z(n14565)
         );
  CND3XL U13703 ( .A(n15274), .B(n14868), .C(entrophy[12]), .Z(n14557) );
  COR2X1 U13704 ( .A(n15349), .B(n14472), .Z(n14936) );
  COND3XL U13705 ( .A(n17808), .B(n15351), .C(n14987), .D(n15060), .Z(n14563)
         );
  CNR2X1 U13706 ( .A(n14559), .B(n14567), .Z(n15197) );
  CANR1X1 U13707 ( .A(datain[2]), .B(n14695), .C(n15197), .Z(n14599) );
  COND3X1 U13708 ( .A(n14561), .B(n14568), .C(n14599), .D(n14560), .Z(n14562)
         );
  CNR2X1 U13709 ( .A(n14969), .B(n14927), .Z(n15198) );
  CANR3XL U13710 ( .A(n15052), .B(n14566), .C(n15198), .D(n14866), .Z(n14569)
         );
  CNR2X2 U13711 ( .A(n14568), .B(n14567), .Z(n14819) );
  CND2XL U13712 ( .A(n14819), .B(dataselector[25]), .Z(n15139) );
  COR2X1 U13713 ( .A(n14559), .B(n14926), .Z(n15064) );
  CND3XL U13714 ( .A(n15139), .B(n14569), .C(n15064), .Z(n14573) );
  CIVX2 U13715 ( .A(n14570), .Z(n14572) );
  CNR4X1 U13716 ( .A(n14573), .B(n15199), .C(n14572), .D(n14571), .Z(n14585)
         );
  CIVX2 U13717 ( .A(n14574), .Z(n14691) );
  CIVX1 U13718 ( .A(n14575), .Z(n14581) );
  COR2XL U13719 ( .A(n14652), .B(n14576), .Z(n14577) );
  CND2XL U13720 ( .A(n15335), .B(n14577), .Z(n14580) );
  CAN8X1 U13721 ( .A(n15064), .B(n14583), .C(n14691), .D(n14582), .E(n14581), 
        .F(n14580), .G(n14579), .H(n14578), .Z(n14584) );
  COR3X1 U13722 ( .A(n14585), .B(n15334), .C(n14584), .Z(n14608) );
  CNR2IX1 U13723 ( .B(entrophy[31]), .A(n17799), .Z(n14586) );
  CNR2X1 U13724 ( .A(n14587), .B(n14586), .Z(n14637) );
  CNR2IX1 U13725 ( .B(n14589), .A(n14588), .Z(n14591) );
  CAN4X1 U13726 ( .A(n14591), .B(n14689), .C(n14590), .D(n15227), .Z(n14592)
         );
  CND2X1 U13727 ( .A(n14819), .B(n15798), .Z(n15081) );
  COND3X1 U13728 ( .A(n14637), .B(n14593), .C(n14592), .D(n15081), .Z(n14594)
         );
  CAN2X1 U13729 ( .A(n14594), .B(n15309), .Z(n14606) );
  CIVX1 U13730 ( .A(n15061), .Z(n14602) );
  CND2X1 U13731 ( .A(n12019), .B(entrophy[22]), .Z(n14597) );
  CNR2X1 U13732 ( .A(n15351), .B(n14966), .Z(n14595) );
  CNR2X1 U13733 ( .A(n14595), .B(n15198), .Z(n14596) );
  CAN3X1 U13734 ( .A(n14597), .B(n14596), .C(n14846), .Z(n14598) );
  CND3XL U13735 ( .A(n14600), .B(n14599), .C(n14598), .Z(n14601) );
  CNR2X1 U13736 ( .A(n14602), .B(n14601), .Z(n14604) );
  CND2XL U13737 ( .A(n15673), .B(scrambler[25]), .Z(n14603) );
  COND1X1 U13738 ( .A(n15112), .B(n14604), .C(n14603), .Z(n14605) );
  CNR2X1 U13739 ( .A(n14606), .B(n14605), .Z(n14607) );
  CND2X1 U13740 ( .A(n14608), .B(n14607), .Z(n8725) );
  COND1XL U13741 ( .A(poly7_shifted[349]), .B(n18228), .C(n18227), .Z(n14610)
         );
  CMXI2X1 U13742 ( .A0(n14610), .A1(n14609), .S(n13040), .Z(n9755) );
  CND2XL U13743 ( .A(n17668), .B(poly7_shifted[379]), .Z(n14612) );
  CND2X1 U13744 ( .A(n12206), .B(poly7_shifted[391]), .Z(n14611) );
  COND4CX1 U13745 ( .A(n14612), .B(n17741), .C(n12206), .D(n14611), .Z(n9725)
         );
  CEOX1 U13746 ( .A(Poly4[51]), .B(n14613), .Z(n14622) );
  CENX1 U13747 ( .A(n14615), .B(n14614), .Z(n14616) );
  CENX1 U13748 ( .A(n14622), .B(n14616), .Z(n14619) );
  COND1XL U13749 ( .A(Poly4[21]), .B(n14619), .C(n17453), .Z(n14618) );
  CMXI2X1 U13750 ( .A0(n14754), .A1(Poly4[38]), .S(n12153), .Z(n14617) );
  COND4CX1 U13751 ( .A(n14619), .B(Poly4[21]), .C(n14618), .D(n14617), .Z(
        n8818) );
  CENX1 U13752 ( .A(Poly4[56]), .B(n14620), .Z(n14621) );
  CENX1 U13753 ( .A(n14622), .B(n14621), .Z(n14625) );
  CIVX2 U13754 ( .A(n15673), .Z(n16435) );
  COND1XL U13755 ( .A(Poly4[35]), .B(n14625), .C(n16435), .Z(n14624) );
  CMXI2X1 U13756 ( .A0(n18082), .A1(Poly4[52]), .S(n12153), .Z(n14623) );
  COND4CX1 U13757 ( .A(n14625), .B(Poly4[35]), .C(n14624), .D(n14623), .Z(
        n8804) );
  COND1XL U13758 ( .A(Poly7[178]), .B(Poly7[399]), .C(n17203), .Z(n14627) );
  CMXI2X1 U13759 ( .A0(n18105), .A1(Poly7[190]), .S(n12977), .Z(n14626) );
  COND4CX1 U13760 ( .A(Poly7[399]), .B(Poly7[178]), .C(n14627), .D(n14626), 
        .Z(n9914) );
  COND1XL U13761 ( .A(Poly7[400]), .B(Poly7[179]), .C(n17449), .Z(n14629) );
  CMXI2X1 U13762 ( .A0(n14436), .A1(Poly7[191]), .S(n12977), .Z(n14628) );
  COND4CX1 U13763 ( .A(Poly7[179]), .B(Poly7[400]), .C(n14629), .D(n14628), 
        .Z(n9913) );
  CNR2X1 U13764 ( .A(n15283), .B(n14850), .Z(n15090) );
  COND11X1 U13765 ( .A(n15090), .B(n14631), .C(n14630), .D(n12216), .Z(n14636)
         );
  CNR2X1 U13766 ( .A(n14652), .B(entrophy[13]), .Z(n14632) );
  CNR3XL U13767 ( .A(n14650), .B(n15798), .C(n14645), .Z(n14634) );
  CANR1XL U13768 ( .A(scrambler[30]), .B(n17959), .C(n14634), .Z(n14635) );
  COND3X1 U13769 ( .A(n14637), .B(n12055), .C(n14636), .D(n14635), .Z(n14679)
         );
  CND2XL U13770 ( .A(n14826), .B(entrophy[22]), .Z(n14639) );
  CANR1X1 U13771 ( .A(datain[5]), .B(n17797), .C(n14819), .Z(n14646) );
  CNR2IX1 U13772 ( .B(n14652), .A(n14646), .Z(n14654) );
  COND1X1 U13773 ( .A(n17809), .B(n15301), .C(n14647), .Z(n14648) );
  CNR3X2 U13774 ( .A(n14648), .B(n17768), .C(n14669), .Z(n14651) );
  CND2XL U13775 ( .A(n15101), .B(datain[0]), .Z(n14649) );
  COND3X1 U13776 ( .A(n14652), .B(n14651), .C(n14650), .D(n14649), .Z(n14653)
         );
  COND1X2 U13777 ( .A(n14654), .B(n14653), .C(n11969), .Z(n14655) );
  CANR1X2 U13778 ( .A(n14656), .B(n14655), .C(n15334), .Z(n14668) );
  CNR2X1 U13779 ( .A(n17763), .B(dataselector[25]), .Z(n14657) );
  CND2X1 U13780 ( .A(n14658), .B(n14657), .Z(n14666) );
  COR3X1 U13781 ( .A(n14936), .B(n14645), .C(n14686), .Z(n14665) );
  CNR3XL U13782 ( .A(n14660), .B(n14645), .C(n14659), .Z(n14663) );
  CNR2IX1 U13783 ( .B(n14661), .A(n15335), .Z(n14662) );
  CNR2X1 U13784 ( .A(n14663), .B(n14662), .Z(n14664) );
  CND3X1 U13785 ( .A(n14666), .B(n14665), .C(n14664), .Z(n14667) );
  CNR2X2 U13786 ( .A(n14668), .B(n14667), .Z(n14676) );
  COND4CXL U13787 ( .A(n14670), .B(entrophy[12]), .C(n14669), .D(n15145), .Z(
        n14671) );
  COND11XL U13788 ( .A(n15352), .B(n14967), .C(n15293), .D(n14671), .Z(n14673)
         );
  CND2X1 U13789 ( .A(n14673), .B(n14672), .Z(n14675) );
  CND3XL U13790 ( .A(n15354), .B(n14868), .C(entrophy[28]), .Z(n14674) );
  CND4X1 U13791 ( .A(n14677), .B(n14676), .C(n14675), .D(n14674), .Z(n14678)
         );
  COR2X1 U13792 ( .A(n14679), .B(n14678), .Z(n8730) );
  CND2X1 U13793 ( .A(n14680), .B(entrophy[13]), .Z(n14836) );
  CND2X1 U13794 ( .A(n14695), .B(entrophy[1]), .Z(n15062) );
  CIVXL U13795 ( .A(n14681), .Z(n14682) );
  CAN8X1 U13796 ( .A(n14685), .B(n15270), .C(n15191), .D(n14684), .E(n14836), 
        .F(n14683), .G(n15062), .H(n14682), .Z(n14711) );
  CNR2X1 U13797 ( .A(n12018), .B(n14686), .Z(n14694) );
  CIVXL U13798 ( .A(n14694), .Z(n14692) );
  CND2XL U13799 ( .A(n14131), .B(datain[3]), .Z(n14688) );
  CND3XL U13800 ( .A(n17792), .B(datain[5]), .C(n14687), .Z(n14820) );
  CND8X1 U13801 ( .A(n14692), .B(n14691), .C(n14690), .D(n14689), .E(n14688), 
        .F(n15136), .G(n14902), .H(n14820), .Z(n14703) );
  CANR2X1 U13802 ( .A(n14694), .B(n14693), .C(entrophy[10]), .D(n11971), .Z(
        n14701) );
  CND2X1 U13803 ( .A(n14695), .B(entrophy[16]), .Z(n15251) );
  CANR2XL U13804 ( .A(n17774), .B(entrophy[12]), .C(scrambler[24]), .D(n17829), 
        .Z(n14699) );
  CND2X1 U13805 ( .A(n17812), .B(datain[0]), .Z(n14698) );
  CND4X1 U13806 ( .A(n14701), .B(n14700), .C(n14699), .D(n14698), .Z(n14702)
         );
  CND2X1 U13807 ( .A(n14705), .B(n14704), .Z(n14708) );
  COND11X1 U13808 ( .A(n14708), .B(n14707), .C(n14706), .D(n15346), .Z(n14709)
         );
  COND3X1 U13809 ( .A(n14711), .B(n12055), .C(n14709), .D(n14710), .Z(n8724)
         );
  CIVX2 U13810 ( .A(n15673), .Z(n16787) );
  COND1XL U13811 ( .A(Poly7[401]), .B(Poly7[180]), .C(n16787), .Z(n14713) );
  CMXI2X1 U13812 ( .A0(n12010), .A1(Poly7[192]), .S(n17273), .Z(n14712) );
  COND4CX1 U13813 ( .A(Poly7[180]), .B(Poly7[401]), .C(n14713), .D(n14712), 
        .Z(n9912) );
  COND1XL U13814 ( .A(Poly7[403]), .B(Poly7[182]), .C(n18234), .Z(n14715) );
  CMXI2X1 U13815 ( .A0(n12415), .A1(Poly7[194]), .S(n17273), .Z(n14714) );
  COND4CX1 U13816 ( .A(Poly7[182]), .B(Poly7[403]), .C(n14715), .D(n14714), 
        .Z(n9910) );
  COND1XL U13817 ( .A(Poly7[402]), .B(Poly7[181]), .C(n17317), .Z(n14718) );
  CMXI2X1 U13818 ( .A0(n14716), .A1(Poly7[193]), .S(n17273), .Z(n14717) );
  COND4CX1 U13819 ( .A(Poly7[181]), .B(Poly7[402]), .C(n14718), .D(n14717), 
        .Z(n9911) );
  CEOXL U13820 ( .A(Poly7[399]), .B(Poly7[183]), .Z(n14721) );
  COND1XL U13821 ( .A(\dataselector_shifted[0] ), .B(n14721), .C(n17298), .Z(
        n14720) );
  CMXI2X1 U13822 ( .A0(n18053), .A1(poly7_shifted[207]), .S(n17273), .Z(n14719) );
  COND4CX1 U13823 ( .A(n14721), .B(\dataselector_shifted[0] ), .C(n14720), .D(
        n14719), .Z(n9909) );
  COND1XL U13824 ( .A(Poly14[210]), .B(Poly14[296]), .C(n17352), .Z(n14723) );
  CMXI2X1 U13825 ( .A0(n13428), .A1(poly14_shifted[242]), .S(n16694), .Z(
        n14722) );
  COND4CX1 U13826 ( .A(Poly14[296]), .B(Poly14[210]), .C(n14723), .D(n14722), 
        .Z(n10179) );
  CIVX2 U13827 ( .A(n15673), .Z(n17375) );
  COND1XL U13828 ( .A(Poly14[300]), .B(Poly14[214]), .C(n17375), .Z(n14725) );
  CMXI2X1 U13829 ( .A0(n14754), .A1(poly14_shifted[246]), .S(n16694), .Z(
        n14724) );
  COND4CX1 U13830 ( .A(Poly14[214]), .B(Poly14[300]), .C(n14725), .D(n14724), 
        .Z(n10175) );
  COND1XL U13831 ( .A(Poly14[297]), .B(Poly14[211]), .C(n17523), .Z(n14727) );
  CMXI2X1 U13832 ( .A0(n18053), .A1(poly14_shifted[243]), .S(n16694), .Z(
        n14726) );
  COND4CX1 U13833 ( .A(Poly14[211]), .B(Poly14[297]), .C(n14727), .D(n14726), 
        .Z(n10178) );
  COND1XL U13834 ( .A(Poly14[295]), .B(Poly14[209]), .C(n17280), .Z(n14729) );
  CIVXL U13835 ( .A(n17711), .Z(n14765) );
  CMXI2X1 U13836 ( .A0(n14765), .A1(poly14_shifted[241]), .S(n16694), .Z(
        n14728) );
  COND4CX1 U13837 ( .A(Poly14[209]), .B(Poly14[295]), .C(n14729), .D(n14728), 
        .Z(n10180) );
  COND1XL U13838 ( .A(Poly14[299]), .B(Poly14[213]), .C(n16372), .Z(n14731) );
  CMXI2X1 U13839 ( .A0(n11996), .A1(poly14_shifted[245]), .S(n16694), .Z(
        n14730) );
  COND4CX1 U13840 ( .A(Poly14[213]), .B(Poly14[299]), .C(n14731), .D(n14730), 
        .Z(n10176) );
  CEOXL U13841 ( .A(Poly14[287]), .B(Poly14[201]), .Z(n14734) );
  COND1XL U13842 ( .A(Poly14[293]), .B(n14734), .C(n18234), .Z(n14733) );
  CMXI2X1 U13843 ( .A0(n18249), .A1(poly14_shifted[233]), .S(n12202), .Z(
        n14732) );
  COND4CX1 U13844 ( .A(n14734), .B(Poly14[293]), .C(n14733), .D(n14732), .Z(
        n10188) );
  COND1XL U13845 ( .A(Poly14[296]), .B(Poly14[176]), .C(n17375), .Z(n14736) );
  CMXI2X1 U13846 ( .A0(n12010), .A1(poly14_shifted[208]), .S(n12202), .Z(
        n14735) );
  COND4CX1 U13847 ( .A(Poly14[176]), .B(Poly14[296]), .C(n14736), .D(n14735), 
        .Z(n10213) );
  COND1XL U13848 ( .A(Poly14[299]), .B(Poly14[179]), .C(n17285), .Z(n14738) );
  CMXI2X1 U13849 ( .A0(n18053), .A1(Poly14[195]), .S(n12202), .Z(n14737) );
  COND4CX1 U13850 ( .A(Poly14[179]), .B(Poly14[299]), .C(n14738), .D(n14737), 
        .Z(n10210) );
  COND1XL U13851 ( .A(Poly14[194]), .B(Poly14[286]), .C(n18234), .Z(n14740) );
  CMXI2X1 U13852 ( .A0(n18210), .A1(Poly14[210]), .S(n12202), .Z(n14739) );
  COND4CX1 U13853 ( .A(Poly14[286]), .B(Poly14[194]), .C(n14740), .D(n14739), 
        .Z(n10195) );
  CEOXL U13854 ( .A(Poly14[296]), .B(Poly14[204]), .Z(n14743) );
  COND1XL U13855 ( .A(Poly14[290]), .B(n14743), .C(n18017), .Z(n14742) );
  COND4CX1 U13856 ( .A(n14743), .B(Poly14[290]), .C(n14742), .D(n14741), .Z(
        n10185) );
  CEOXL U13857 ( .A(Poly14[286]), .B(Poly14[200]), .Z(n14746) );
  COND1XL U13858 ( .A(Poly14[292]), .B(n14746), .C(n17998), .Z(n14745) );
  CMXI2X1 U13859 ( .A0(n13994), .A1(poly14_shifted[232]), .S(n12202), .Z(
        n14744) );
  COND4CX1 U13860 ( .A(n14746), .B(Poly14[292]), .C(n14745), .D(n14744), .Z(
        n10189) );
  COND1XL U13861 ( .A(Poly14[285]), .B(Poly14[193]), .C(n17453), .Z(n14748) );
  CMXI2X1 U13862 ( .A0(n18048), .A1(Poly14[209]), .S(n12202), .Z(n14747) );
  COND4CX1 U13863 ( .A(Poly14[193]), .B(Poly14[285]), .C(n14748), .D(n14747), 
        .Z(n10196) );
  CEOXL U13864 ( .A(Poly14[299]), .B(Poly14[207]), .Z(n14751) );
  COND1XL U13865 ( .A(Poly14[293]), .B(n14751), .C(n18047), .Z(n14750) );
  CMXI2X1 U13866 ( .A0(n12003), .A1(poly14_shifted[239]), .S(n12202), .Z(
        n14749) );
  COND4CX1 U13867 ( .A(n14751), .B(Poly14[293]), .C(n14750), .D(n14749), .Z(
        n10182) );
  COND1XL U13868 ( .A(Poly14[298]), .B(Poly14[178]), .C(n17285), .Z(n14753) );
  CMXI2X1 U13869 ( .A0(n12415), .A1(Poly14[194]), .S(n12202), .Z(n14752) );
  COND4CX1 U13870 ( .A(Poly14[178]), .B(Poly14[298]), .C(n14753), .D(n14752), 
        .Z(n10211) );
  COND1XL U13871 ( .A(Poly7[409]), .B(Poly7[58]), .C(n17538), .Z(n14756) );
  CMXI2X1 U13872 ( .A0(n14754), .A1(poly7_shifted[82]), .S(n17471), .Z(n14755)
         );
  COND4CX1 U13873 ( .A(Poly7[58]), .B(Poly7[409]), .C(n14756), .D(n14755), .Z(
        n10034) );
  CIVX2 U13874 ( .A(n15673), .Z(n17458) );
  COND1XL U13875 ( .A(Poly7[405]), .B(Poly7[54]), .C(n17458), .Z(n14758) );
  CMXI2X1 U13876 ( .A0(n13428), .A1(poly7_shifted[78]), .S(n17471), .Z(n14757)
         );
  COND4CX1 U13877 ( .A(Poly7[54]), .B(Poly7[405]), .C(n14758), .D(n14757), .Z(
        n10038) );
  COND1XL U13878 ( .A(Poly7[403]), .B(Poly7[52]), .C(n17453), .Z(n14760) );
  CMXI2X1 U13879 ( .A0(n12010), .A1(poly7_shifted[76]), .S(n17471), .Z(n14759)
         );
  COND4CX1 U13880 ( .A(Poly7[52]), .B(Poly7[403]), .C(n14760), .D(n14759), .Z(
        n10040) );
  COND1XL U13881 ( .A(Poly7[406]), .B(Poly7[55]), .C(n17398), .Z(n14762) );
  CMXI2X1 U13882 ( .A0(n18053), .A1(poly7_shifted[79]), .S(n17471), .Z(n14761)
         );
  COND4CX1 U13883 ( .A(Poly7[55]), .B(Poly7[406]), .C(n14762), .D(n14761), .Z(
        n10037) );
  COND1XL U13884 ( .A(Poly7[407]), .B(Poly7[56]), .C(n17538), .Z(n14764) );
  CMXI2X1 U13885 ( .A0(n12004), .A1(poly7_shifted[80]), .S(n17471), .Z(n14763)
         );
  COND4CX1 U13886 ( .A(Poly7[56]), .B(Poly7[407]), .C(n14764), .D(n14763), .Z(
        n10036) );
  COND1XL U13887 ( .A(\dataselector_shifted[0] ), .B(Poly7[53]), .C(n17063), 
        .Z(n14767) );
  CMXI2X1 U13888 ( .A0(n14765), .A1(poly7_shifted[77]), .S(n17471), .Z(n14766)
         );
  COND4CX1 U13889 ( .A(Poly7[53]), .B(\dataselector_shifted[0] ), .C(n14767), 
        .D(n14766), .Z(n10039) );
  COND1XL U13890 ( .A(Poly7[408]), .B(Poly7[57]), .C(n17362), .Z(n14769) );
  CMXI2X1 U13891 ( .A0(n11988), .A1(poly7_shifted[81]), .S(n17471), .Z(n14768)
         );
  COND4CX1 U13892 ( .A(Poly7[57]), .B(Poly7[408]), .C(n14769), .D(n14768), .Z(
        n10035) );
  COND1XL U13893 ( .A(Poly7[410]), .B(Poly7[59]), .C(n17705), .Z(n14771) );
  CMXI2X1 U13894 ( .A0(n18138), .A1(poly7_shifted[83]), .S(n17471), .Z(n14770)
         );
  COND4CX1 U13895 ( .A(Poly7[59]), .B(Poly7[410]), .C(n14771), .D(n14770), .Z(
        n10033) );
  CANR4CX1 U13896 ( .A(Poly2[38]), .B(n14772), .C(n17571), .D(n17306), .Z(
        n14775) );
  CANR2X1 U13897 ( .A(n17306), .B(Poly2[50]), .C(n14773), .D(Poly2[38]), .Z(
        n14774) );
  CND2IX1 U13898 ( .B(n14775), .A(n14774), .Z(n8960) );
  COND1XL U13899 ( .A(Poly4[17]), .B(n14778), .C(n17598), .Z(n14777) );
  CMXI2X1 U13900 ( .A0(n13428), .A1(Poly4[34]), .S(n12153), .Z(n14776) );
  COND4CX1 U13901 ( .A(n14778), .B(Poly4[17]), .C(n14777), .D(n14776), .Z(
        n8822) );
  CANR2X1 U13902 ( .A(n17775), .B(datain[2]), .C(datain[4]), .D(n17774), .Z(
        n14787) );
  CANR2X1 U13903 ( .A(n17812), .B(entrophy[1]), .C(entrophy[24]), .D(n11971), 
        .Z(n14786) );
  CIVX2 U13904 ( .A(n14779), .Z(n15007) );
  CANR2XL U13905 ( .A(n15007), .B(n15314), .C(scrambler[13]), .D(n17826), .Z(
        n14785) );
  CND2XL U13906 ( .A(n15052), .B(datain[0]), .Z(n14780) );
  COND3X1 U13907 ( .A(n15229), .B(n14928), .C(n14781), .D(n14780), .Z(n14783)
         );
  CND3XL U13908 ( .A(n14783), .B(n12216), .C(n14782), .Z(n14784) );
  CAN4X1 U13909 ( .A(n14787), .B(n14786), .C(n14785), .D(n14784), .Z(n14816)
         );
  COND1XL U13910 ( .A(n15052), .B(entrophy[16]), .C(n15034), .Z(n14793) );
  CND2X1 U13911 ( .A(n15354), .B(entrophy[14]), .Z(n15103) );
  CIVX1 U13912 ( .A(n15103), .Z(n14791) );
  CND2XL U13913 ( .A(n11969), .B(n17805), .Z(n14789) );
  CNR3XL U13914 ( .A(n14789), .B(n14788), .C(n14795), .Z(n14790) );
  CANR3X1 U13915 ( .A(n14864), .B(n17792), .C(n14791), .D(n14790), .Z(n14792)
         );
  COND4CX1 U13916 ( .A(n14979), .B(n15211), .C(n14793), .D(n14792), .Z(n14794)
         );
  CND2X1 U13917 ( .A(n17804), .B(n14794), .Z(n14806) );
  CNR2X1 U13918 ( .A(n14969), .B(n14795), .Z(n14800) );
  CNR2XL U13919 ( .A(n14796), .B(n14999), .Z(n14798) );
  CNR2IX1 U13920 ( .B(n14798), .A(n14797), .Z(n14799) );
  CNR2X1 U13921 ( .A(n14800), .B(n14799), .Z(n14801) );
  CND3X1 U13922 ( .A(n14912), .B(n14802), .C(n14801), .Z(n14804) );
  COND11X2 U13923 ( .A(n14804), .B(n14803), .C(n15144), .D(n15346), .Z(n14805)
         );
  CND2X2 U13924 ( .A(n14806), .B(n14805), .Z(n14814) );
  CNR2X1 U13925 ( .A(n13958), .B(n14807), .Z(n15216) );
  CNR2X1 U13926 ( .A(n15218), .B(n14807), .Z(n17790) );
  CNR2X1 U13927 ( .A(n15283), .B(n14808), .Z(n17777) );
  CNR2XL U13928 ( .A(n14226), .B(n14850), .Z(n14810) );
  CNR2X1 U13929 ( .A(n12018), .B(n15352), .Z(n14809) );
  CNR8X1 U13930 ( .A(n15058), .B(n15216), .C(n14811), .D(n17790), .E(n15017), 
        .F(n17777), .G(n14810), .H(n14809), .Z(n14812) );
  CNR2X1 U13931 ( .A(n14812), .B(n15112), .Z(n14813) );
  CNR2X2 U13932 ( .A(n14814), .B(n14813), .Z(n14815) );
  CND2X1 U13933 ( .A(n14816), .B(n14815), .Z(n8713) );
  COND1XL U13934 ( .A(Poly7[410]), .B(Poly7[244]), .C(n16427), .Z(n14818) );
  CMXI2X1 U13935 ( .A0(n12010), .A1(poly7_shifted[268]), .S(n12625), .Z(n14817) );
  COND4CX1 U13936 ( .A(Poly7[244]), .B(Poly7[410]), .C(n14818), .D(n14817), 
        .Z(n9848) );
  CIVXL U13937 ( .A(n14819), .Z(n14821) );
  CND2X1 U13938 ( .A(n14848), .B(entrophy[17]), .Z(n14915) );
  CND3XL U13939 ( .A(n14821), .B(n14915), .C(n14820), .Z(n14822) );
  COND4CX1 U13940 ( .A(entrophy[25]), .B(n15348), .C(n14822), .D(n12216), .Z(
        n14835) );
  CIVX2 U13941 ( .A(n14823), .Z(n14825) );
  CND4X1 U13942 ( .A(n14825), .B(n15257), .C(n14824), .D(n14891), .Z(n14830)
         );
  COND1X1 U13943 ( .A(n14826), .B(n12019), .C(entrophy[15]), .Z(n14828) );
  CND2X1 U13944 ( .A(n15256), .B(entrophy[24]), .Z(n14948) );
  CND3X1 U13945 ( .A(n14828), .B(n14948), .C(n14827), .Z(n14829) );
  COR2X1 U13946 ( .A(n14830), .B(n14829), .Z(n14832) );
  CNR2X1 U13947 ( .A(n15338), .B(n14927), .Z(n14831) );
  CANR1X1 U13948 ( .A(n15346), .B(n14832), .C(n14831), .Z(n14834) );
  CANR2XL U13949 ( .A(n17787), .B(entrophy[22]), .C(scrambler[9]), .D(n17959), 
        .Z(n14833) );
  CND3XL U13950 ( .A(n14835), .B(n14834), .C(n14833), .Z(n14844) );
  CND4X1 U13951 ( .A(n14965), .B(n14837), .C(n14836), .D(n15172), .Z(n14840)
         );
  CND2X1 U13952 ( .A(n14695), .B(entrophy[11]), .Z(n15322) );
  COND1XL U13953 ( .A(dataselector[21]), .B(n15124), .C(n15322), .Z(n15225) );
  CIVX2 U13954 ( .A(n17793), .Z(n14839) );
  CNR4X1 U13955 ( .A(n14840), .B(n15225), .C(n14839), .D(n14838), .Z(n14842)
         );
  CNR2IXL U13956 ( .B(n16249), .A(n14852), .Z(n14841) );
  CNIVX1 U13957 ( .A(n14841), .Z(n15273) );
  CND2X1 U13958 ( .A(n15273), .B(n14866), .Z(n15261) );
  CNR2X1 U13959 ( .A(n14842), .B(n15261), .Z(n14843) );
  CNR2X1 U13960 ( .A(n14844), .B(n14843), .Z(n14856) );
  CND4X1 U13961 ( .A(n15137), .B(n14847), .C(n14846), .D(n14845), .Z(n14854)
         );
  CND2X1 U13962 ( .A(n11974), .B(datain[2]), .Z(n14900) );
  CND2XL U13963 ( .A(n14848), .B(entrophy[20]), .Z(n14849) );
  COND3X1 U13964 ( .A(n14851), .B(n14850), .C(n14900), .D(n14849), .Z(n14853)
         );
  CNR3XL U13965 ( .A(n14852), .B(n16249), .C(n14866), .Z(n15288) );
  COND1XL U13966 ( .A(n14854), .B(n14853), .C(n15288), .Z(n14855) );
  CND2X1 U13967 ( .A(n14856), .B(n14855), .Z(n8709) );
  CND2X1 U13968 ( .A(n14857), .B(datain[7]), .Z(n14949) );
  CND2XL U13969 ( .A(n15111), .B(entrophy[27]), .Z(n14858) );
  CND4X1 U13970 ( .A(n14860), .B(n14949), .C(n14859), .D(n14858), .Z(n14874)
         );
  CND3XL U13971 ( .A(n15274), .B(n14868), .C(entrophy[13]), .Z(n14863) );
  CNR2IX1 U13972 ( .B(entrophy[20]), .A(n14958), .Z(n14861) );
  COND3X1 U13973 ( .A(n11970), .B(n15339), .C(n14863), .D(n14862), .Z(n14873)
         );
  CIVX1 U13974 ( .A(n17787), .Z(n15107) );
  CIVXL U13975 ( .A(n14864), .Z(n14865) );
  CANR4CX1 U13976 ( .A(n14866), .B(n14226), .C(n14865), .D(n14645), .Z(n14867)
         );
  COND4CX1 U13977 ( .A(datain[6]), .B(n14913), .C(n17770), .D(n14867), .Z(
        n14870) );
  CND3XL U13978 ( .A(n14976), .B(entrophy[7]), .C(n14868), .Z(n14869) );
  COND3X1 U13979 ( .A(n15107), .B(n14871), .C(n14870), .D(n14869), .Z(n14872)
         );
  CANR3X1 U13980 ( .A(n15145), .B(n14874), .C(n14873), .D(n14872), .Z(n14899)
         );
  CND2XL U13981 ( .A(n14875), .B(entrophy[17]), .Z(n14876) );
  CANR1XL U13982 ( .A(n14936), .B(n14979), .C(n14876), .Z(n14885) );
  CANR2XL U13983 ( .A(n14878), .B(n14877), .C(scrambler[19]), .D(n17744), .Z(
        n14882) );
  CND3XL U13984 ( .A(n14880), .B(n14868), .C(n14879), .Z(n14881) );
  COND3X1 U13985 ( .A(n14883), .B(n17800), .C(n14882), .D(n14881), .Z(n14884)
         );
  CND3XL U13986 ( .A(n14892), .B(n14891), .C(n14890), .Z(n14897) );
  COND3X1 U13987 ( .A(n14895), .B(n14894), .C(n14893), .D(n14988), .Z(n14896)
         );
  COND1XL U13988 ( .A(n14897), .B(n14896), .C(n15220), .Z(n14898) );
  CND2XL U13989 ( .A(n14695), .B(entrophy[27]), .Z(n14903) );
  CAN8X1 U13990 ( .A(n14905), .B(n15268), .C(n14904), .D(n14903), .E(n14902), 
        .F(n14901), .G(n14900), .H(n15217), .Z(n14942) );
  CND2XL U13991 ( .A(n15034), .B(entrophy[22]), .Z(n14907) );
  CND2XL U13992 ( .A(n17767), .B(entrophy[16]), .Z(n14906) );
  CMXI2X1 U13993 ( .A0(n14907), .A1(n14906), .S(n14928), .Z(n14923) );
  CND2X1 U13994 ( .A(n15043), .B(entrophy[9]), .Z(n15153) );
  CND2X1 U13995 ( .A(n17812), .B(entrophy[7]), .Z(n14911) );
  COND2X1 U13996 ( .A(n17778), .B(n14909), .C(n15108), .D(n17784), .Z(n14910)
         );
  CNR2IX1 U13997 ( .B(n14911), .A(n14910), .Z(n14920) );
  CND2X1 U13998 ( .A(n14912), .B(n15025), .Z(n14918) );
  CANR2X1 U13999 ( .A(n14913), .B(entrophy[27]), .C(entrophy[1]), .D(n15052), 
        .Z(n14914) );
  CND2X1 U14000 ( .A(n14915), .B(n14914), .Z(n14916) );
  CANR2X1 U14001 ( .A(n14918), .B(n14917), .C(n15145), .D(n14916), .Z(n14919)
         );
  CND3X2 U14002 ( .A(n14921), .B(n14920), .C(n14919), .Z(n14922) );
  CANR1X1 U14003 ( .A(n14923), .B(n17804), .C(n14922), .Z(n14941) );
  COND3XL U14004 ( .A(n15218), .B(n14926), .C(n14925), .D(n14924), .Z(n14939)
         );
  CNR4X1 U14005 ( .A(n14928), .B(n17799), .C(n12055), .D(n14927), .Z(n14929)
         );
  CANR1XL U14006 ( .A(scrambler[11]), .B(n17744), .C(n14929), .Z(n14932) );
  COR2X1 U14007 ( .A(n14930), .B(n15335), .Z(n14931) );
  CND2X1 U14008 ( .A(n14932), .B(n14931), .Z(n14938) );
  COND4CX1 U14009 ( .A(n14936), .B(n14935), .C(n14934), .D(n14933), .Z(n14937)
         );
  COND3X1 U14010 ( .A(n14942), .B(n15236), .C(n14941), .D(n14940), .Z(n8711)
         );
  CEOXL U14011 ( .A(n14943), .B(dataselector[12]), .Z(n14945) );
  COND2XL U14012 ( .A(n14945), .B(n17959), .C(n17654), .D(n14944), .Z(n14946)
         );
  CAOR1X1 U14013 ( .A(n16410), .B(dataselector[19]), .C(n14946), .Z(n8776) );
  CAN4X1 U14014 ( .A(n15227), .B(n14949), .C(n14948), .D(n14947), .Z(n14954)
         );
  CANR2X1 U14015 ( .A(n17787), .B(entrophy[13]), .C(scrambler[4]), .D(n17259), 
        .Z(n14953) );
  CANR2X1 U14016 ( .A(n17770), .B(n14951), .C(n15346), .D(n14950), .Z(n14952)
         );
  COND3X1 U14017 ( .A(n14954), .B(n15170), .C(n14953), .D(n14952), .Z(n14997)
         );
  COND11X1 U14018 ( .A(n14957), .B(n14956), .C(n14955), .D(n15220), .Z(n14995)
         );
  CNR2IXL U14019 ( .B(entrophy[1]), .A(n14958), .Z(n14959) );
  CAN2X1 U14020 ( .A(n15256), .B(entrophy[12]), .Z(n15065) );
  CIVXL U14021 ( .A(n14960), .Z(n14961) );
  CNR3X2 U14022 ( .A(n15065), .B(n14962), .C(n14961), .Z(n14964) );
  CANR11X1 U14023 ( .A(n14965), .B(n15097), .C(n14964), .D(n14963), .Z(n14974)
         );
  CANR2X1 U14024 ( .A(n14969), .B(n14968), .C(n14967), .D(n14966), .Z(n14971)
         );
  CANR2X1 U14025 ( .A(datain[7]), .B(n15074), .C(n14971), .D(n14970), .Z(
        n14972) );
  CNR2X1 U14026 ( .A(n14972), .B(n17785), .Z(n14973) );
  CNR3X1 U14027 ( .A(n14975), .B(n14974), .C(n14973), .Z(n14994) );
  CANR2X1 U14028 ( .A(n15354), .B(entrophy[26]), .C(entrophy[3]), .D(n14976), 
        .Z(n14978) );
  CANR4CX1 U14029 ( .A(n15219), .B(n14979), .C(n14978), .D(n14645), .Z(n14980)
         );
  CIVX2 U14030 ( .A(n14980), .Z(n14993) );
  CNR2XL U14031 ( .A(n14981), .B(n15106), .Z(n14984) );
  CNR2X1 U14032 ( .A(n15005), .B(n14982), .Z(n14983) );
  CND2IX1 U14033 ( .B(n14984), .A(n14983), .Z(n14991) );
  CIVXL U14034 ( .A(n14985), .Z(n14989) );
  CAN4X1 U14035 ( .A(n14995), .B(n14994), .C(n14993), .D(n14992), .Z(n14996)
         );
  CND2IX1 U14036 ( .B(n14997), .A(n14996), .Z(n8704) );
  CIVXL U14037 ( .A(n14998), .Z(n15004) );
  CNR2X1 U14038 ( .A(n15283), .B(n14999), .Z(n15192) );
  CANR1XL U14039 ( .A(datain[6]), .B(n14695), .C(n15192), .Z(n15000) );
  CND2X1 U14040 ( .A(n15206), .B(entrophy[14]), .Z(n15258) );
  COND3XL U14041 ( .A(n15001), .B(n15218), .C(n15000), .D(n15258), .Z(n15002)
         );
  COR4X1 U14042 ( .A(n15295), .B(n15004), .C(n15003), .D(n15002), .Z(n15016)
         );
  COR3X1 U14043 ( .A(n15007), .B(n15006), .C(n15005), .Z(n15011) );
  CND2X1 U14044 ( .A(n15009), .B(n15008), .Z(n15010) );
  CNR2X1 U14045 ( .A(n15011), .B(n15010), .Z(n15014) );
  CANR2XL U14046 ( .A(n17787), .B(datain[5]), .C(scrambler[7]), .D(n17495), 
        .Z(n15013) );
  CANR2X1 U14047 ( .A(n17812), .B(entrophy[27]), .C(entrophy[7]), .D(n17774), 
        .Z(n15012) );
  COND3X1 U14048 ( .A(n15014), .B(n17778), .C(n15013), .D(n15012), .Z(n15015)
         );
  CANR1X1 U14049 ( .A(n15220), .B(n15016), .C(n15015), .Z(n15032) );
  CIVXL U14050 ( .A(n15141), .Z(n15019) );
  CNR2X1 U14051 ( .A(n14226), .B(n15044), .Z(n15212) );
  COR8X1 U14052 ( .A(n15021), .B(n15020), .C(n15019), .D(n15018), .E(n15212), 
        .F(n15091), .G(n17790), .H(n15017), .Z(n15030) );
  CND2X1 U14053 ( .A(n13945), .B(entrophy[13]), .Z(n15134) );
  CIVX1 U14054 ( .A(n15022), .Z(n15027) );
  CND2X1 U14055 ( .A(n11974), .B(entrophy[22]), .Z(n15343) );
  CIVX1 U14056 ( .A(n15023), .Z(n15026) );
  CND8X1 U14057 ( .A(n15134), .B(n15064), .C(n15028), .D(n15027), .E(n15343), 
        .F(n15026), .G(n15025), .H(n15024), .Z(n15029) );
  CANR2X1 U14058 ( .A(n15030), .B(n15309), .C(n15145), .D(n15029), .Z(n15031)
         );
  CND2X1 U14059 ( .A(n15032), .B(n15031), .Z(n8707) );
  CIVXL U14060 ( .A(scrambler[20]), .Z(n15038) );
  CND2X1 U14061 ( .A(n15034), .B(n15033), .Z(n15037) );
  CND3XL U14062 ( .A(n12216), .B(n15035), .C(entrophy[26]), .Z(n15036) );
  COND3XL U14063 ( .A(n12031), .B(n15038), .C(n15037), .D(n15036), .Z(n15039)
         );
  CANR1XL U14064 ( .A(entrophy[6]), .B(n17774), .C(n15039), .Z(n15040) );
  COAN1X1 U14065 ( .A(n15334), .B(n15041), .C(n15040), .Z(n15086) );
  CNR2XL U14066 ( .A(n15042), .B(n15175), .Z(n15158) );
  CANR2XL U14067 ( .A(n15043), .B(n15158), .C(datain[6]), .D(n17812), .Z(
        n15057) );
  COR3X1 U14068 ( .A(n15168), .B(n15044), .C(n15334), .Z(n15056) );
  CIVXL U14069 ( .A(n15047), .Z(n15048) );
  CANR1X1 U14070 ( .A(n15251), .B(n15329), .C(n15048), .Z(n15049) );
  CANR1X1 U14071 ( .A(entrophy[3]), .B(n17787), .C(n15049), .Z(n15050) );
  CND2X1 U14072 ( .A(n15052), .B(datain[2]), .Z(n17801) );
  COR2XL U14073 ( .A(n17801), .B(dataselector[25]), .Z(n15054) );
  CND3X1 U14074 ( .A(n15057), .B(n15056), .C(n15055), .Z(n15084) );
  CIVX1 U14075 ( .A(n15058), .Z(n15069) );
  CND4X1 U14076 ( .A(n15064), .B(n15063), .C(n15062), .D(n15061), .Z(n15066)
         );
  CNR3X1 U14077 ( .A(n15067), .B(n15066), .C(n15065), .Z(n15068) );
  CANR1X1 U14078 ( .A(n15069), .B(n15068), .C(n15236), .Z(n15083) );
  CND2XL U14079 ( .A(n15071), .B(n15070), .Z(n15073) );
  CANR3X1 U14080 ( .A(n15074), .B(entrophy[31]), .C(n15073), .D(n15072), .Z(
        n15080) );
  COND1XL U14081 ( .A(n15339), .B(n15076), .C(n15075), .Z(n15078) );
  CND2XL U14082 ( .A(n15168), .B(n17808), .Z(n15077) );
  CND2X1 U14083 ( .A(n15078), .B(n15077), .Z(n15079) );
  CANR11X1 U14084 ( .A(n15081), .B(n15080), .C(n15079), .D(n15112), .Z(n15082)
         );
  CNR3X2 U14085 ( .A(n15084), .B(n15083), .C(n15082), .Z(n15085) );
  CND2X1 U14086 ( .A(n15086), .B(n15085), .Z(n8720) );
  CENX1 U14087 ( .A(Poly4[54]), .B(n15640), .Z(n15087) );
  CENX1 U14088 ( .A(n17326), .B(n15087), .Z(n15183) );
  CIVX2 U14089 ( .A(n15673), .Z(n16307) );
  COND1XL U14090 ( .A(Poly4[26]), .B(n15183), .C(n16307), .Z(n15089) );
  CMXI2X1 U14091 ( .A0(n16381), .A1(Poly4[43]), .S(n12153), .Z(n15088) );
  COND4CX1 U14092 ( .A(n15183), .B(Poly4[26]), .C(n15089), .D(n15088), .Z(
        n8813) );
  CIVX2 U14093 ( .A(n15090), .Z(n15350) );
  CIVXL U14094 ( .A(n15091), .Z(n15092) );
  CAN8X1 U14095 ( .A(n15097), .B(n15350), .C(n15096), .D(n15095), .E(n15268), 
        .F(n15094), .G(n15093), .H(n15092), .Z(n15129) );
  CIVXL U14096 ( .A(n15098), .Z(n15100) );
  CANR1XL U14097 ( .A(n15101), .B(n15100), .C(n15099), .Z(n15102) );
  COND3X1 U14098 ( .A(n15104), .B(n17808), .C(n15103), .D(n15102), .Z(n15118)
         );
  CANR2X1 U14099 ( .A(n15309), .B(n15313), .C(scrambler[27]), .D(n17495), .Z(
        n15105) );
  COND4CX1 U14100 ( .A(n15108), .B(n15107), .C(n15106), .D(n15105), .Z(n15117)
         );
  CANR2XL U14101 ( .A(n15111), .B(entrophy[16]), .C(n15110), .D(n15109), .Z(
        n15113) );
  CANR11X1 U14102 ( .A(n15115), .B(n15114), .C(n15113), .D(n15112), .Z(n15116)
         );
  CANR3X1 U14103 ( .A(n14868), .B(n15118), .C(n15117), .D(n15116), .Z(n15128)
         );
  CAN2XL U14104 ( .A(n15119), .B(entrophy[14]), .Z(n15122) );
  CND2X1 U14105 ( .A(n17759), .B(entrophy[23]), .Z(n15132) );
  CND3XL U14106 ( .A(n15141), .B(n15120), .C(n15132), .Z(n15121) );
  COR2X1 U14107 ( .A(n15122), .B(n15121), .Z(n15126) );
  CANR2X1 U14108 ( .A(entrophy[24]), .B(n15330), .C(entrophy[13]), .D(n11971), 
        .Z(n15123) );
  COND4CX1 U14109 ( .A(n15124), .B(n17794), .C(n17800), .D(n15123), .Z(n15125)
         );
  CANR1X1 U14110 ( .A(n12216), .B(n15126), .C(n15125), .Z(n15127) );
  COND3X1 U14111 ( .A(n15129), .B(n12055), .C(n15128), .D(n15127), .Z(n8727)
         );
  CIVX1 U14112 ( .A(n15130), .Z(n15135) );
  CIVX1 U14113 ( .A(n15131), .Z(n15133) );
  CAN8X1 U14114 ( .A(n15139), .B(n15138), .C(n15137), .D(n15136), .E(n15135), 
        .F(n15134), .G(n15133), .H(n15132), .Z(n15180) );
  COND3X1 U14115 ( .A(n15211), .B(n15149), .C(n15141), .D(n15140), .Z(n15147)
         );
  COND1XL U14116 ( .A(n15147), .B(n15146), .C(n15145), .Z(n15179) );
  CND3XL U14117 ( .A(n15274), .B(n17804), .C(entrophy[20]), .Z(n15156) );
  COND2XL U14118 ( .A(n15300), .B(n15149), .C(n17799), .D(n15148), .Z(n15152)
         );
  CIVXL U14119 ( .A(n15150), .Z(n15151) );
  COND1XL U14120 ( .A(n15152), .B(n15151), .C(n15220), .Z(n15155) );
  CND3XL U14121 ( .A(n15156), .B(n15155), .C(n15154), .Z(n15177) );
  CND2XL U14122 ( .A(n17770), .B(n15157), .Z(n15167) );
  CND3XL U14123 ( .A(n17792), .B(n17767), .C(n15158), .Z(n15166) );
  COND4CX1 U14124 ( .A(n15160), .B(n11969), .C(n15159), .D(n12216), .Z(n15161)
         );
  CIVX2 U14125 ( .A(n15161), .Z(n15164) );
  CIVXL U14126 ( .A(scrambler[17]), .Z(n15162) );
  CNR2XL U14127 ( .A(n16947), .B(n15162), .Z(n15163) );
  CNR2X1 U14128 ( .A(n15164), .B(n15163), .Z(n15165) );
  CAOR1X1 U14129 ( .A(n15172), .B(n15171), .C(n15170), .Z(n15173) );
  COND3X1 U14130 ( .A(n15230), .B(n15175), .C(n15174), .D(n15173), .Z(n15176)
         );
  CNR2X1 U14131 ( .A(n15177), .B(n15176), .Z(n15178) );
  COND3X1 U14132 ( .A(n15180), .B(n17785), .C(n15179), .D(n15178), .Z(n8717)
         );
  CIVX2 U14133 ( .A(n15673), .Z(n17527) );
  COND1XL U14134 ( .A(Poly4[40]), .B(n15183), .C(n17527), .Z(n15182) );
  CMXI2X1 U14135 ( .A0(n18249), .A1(Poly4[57]), .S(n12153), .Z(n15181) );
  COND4CX1 U14136 ( .A(n15183), .B(Poly4[40]), .C(n15182), .D(n15181), .Z(
        n8799) );
  CND2X1 U14137 ( .A(n17935), .B(poly5_shifted[72]), .Z(n15185) );
  CND2X1 U14138 ( .A(n16787), .B(poly5_shifted[58]), .Z(n15184) );
  COND3X1 U14139 ( .A(n17935), .B(n17735), .C(n15185), .D(n15184), .Z(n11468)
         );
  CENX1 U14140 ( .A(n15187), .B(n15186), .Z(n15245) );
  COND1XL U14141 ( .A(Poly4[38]), .B(n15245), .C(n16323), .Z(n15189) );
  CMXI2X1 U14142 ( .A0(n11999), .A1(Poly4[55]), .S(n12153), .Z(n15188) );
  COND4CX1 U14143 ( .A(n15245), .B(Poly4[38]), .C(n15189), .D(n15188), .Z(
        n8801) );
  CIVX1 U14144 ( .A(n15190), .Z(n15196) );
  CIVX1 U14145 ( .A(n15191), .Z(n15194) );
  CNR8X1 U14146 ( .A(n15199), .B(n15198), .C(n15197), .D(n15196), .E(n15195), 
        .F(n15194), .G(n15193), .H(n15192), .Z(n15237) );
  CNR2X1 U14147 ( .A(n12459), .B(n15333), .Z(n15310) );
  CIVX2 U14148 ( .A(n15310), .Z(n15201) );
  CND2X1 U14149 ( .A(n15202), .B(n15201), .Z(n15204) );
  COR2X1 U14150 ( .A(n15204), .B(n15203), .Z(n15210) );
  CIVXL U14151 ( .A(n15205), .Z(n15207) );
  CND2X1 U14152 ( .A(n14695), .B(entrophy[3]), .Z(n15282) );
  CND2X1 U14153 ( .A(n15206), .B(entrophy[18]), .Z(n15321) );
  CND4X1 U14154 ( .A(n15208), .B(n15207), .C(n15282), .D(n15321), .Z(n15209)
         );
  COND1X1 U14155 ( .A(n15210), .B(n15209), .C(n15145), .Z(n15224) );
  CND2IX1 U14156 ( .B(n15211), .A(n15249), .Z(n15215) );
  CNR2X1 U14157 ( .A(n15213), .B(n15212), .Z(n15214) );
  COND1XL U14158 ( .A(n15219), .B(n15218), .C(n17760), .Z(n15221) );
  COND1X2 U14159 ( .A(n15222), .B(n15221), .C(n15220), .Z(n15223) );
  CAN2X1 U14160 ( .A(n15224), .B(n15223), .Z(n15235) );
  CIVXL U14161 ( .A(n15225), .Z(n15228) );
  CND4X1 U14162 ( .A(n15228), .B(n15227), .C(n17761), .D(n15226), .Z(n15233)
         );
  COND2X1 U14163 ( .A(n15339), .B(n15230), .C(n15338), .D(n15229), .Z(n15232)
         );
  CAOR2XL U14164 ( .A(scrambler[10]), .B(n17829), .C(n17787), .D(datain[6]), 
        .Z(n15231) );
  CANR3X1 U14165 ( .A(n12216), .B(n15233), .C(n15232), .D(n15231), .Z(n15234)
         );
  COND3X1 U14166 ( .A(n15237), .B(n15236), .C(n15235), .D(n15234), .Z(n8710)
         );
  CEOX1 U14167 ( .A(Poly4[50]), .B(Poly4[52]), .Z(n17328) );
  CENX1 U14168 ( .A(n15238), .B(Poly4[36]), .Z(n15239) );
  CENX1 U14169 ( .A(n17328), .B(n15239), .Z(n15242) );
  COND1XL U14170 ( .A(n15651), .B(n15242), .C(n16787), .Z(n15241) );
  CMXI2X1 U14171 ( .A0(n18241), .A1(Poly4[53]), .S(n12153), .Z(n15240) );
  COND4CX1 U14172 ( .A(n15242), .B(n15651), .C(n15241), .D(n15240), .Z(n8803)
         );
  COND1XL U14173 ( .A(n15245), .B(Poly4[24]), .C(n17398), .Z(n15244) );
  CMXI2XL U14174 ( .A0(n12001), .A1(Poly4[41]), .S(n12153), .Z(n15243) );
  COND4CX1 U14175 ( .A(Poly4[24]), .B(n15245), .C(n15244), .D(n15243), .Z(
        n8815) );
  CANR1XL U14176 ( .A(datain[7]), .B(n17759), .C(n15250), .Z(n15253) );
  CAN4X1 U14177 ( .A(n15254), .B(n15253), .C(n15252), .D(n15251), .Z(n15294)
         );
  CANR1X1 U14178 ( .A(entrophy[20]), .B(n15256), .C(n15255), .Z(n15259) );
  CND4X1 U14179 ( .A(n15260), .B(n15259), .C(n15258), .D(n15257), .Z(n15264)
         );
  CIVX1 U14180 ( .A(n15261), .Z(n15262) );
  COND1XL U14181 ( .A(n15264), .B(n15263), .C(n15262), .Z(n15281) );
  CND2X1 U14182 ( .A(n11971), .B(entrophy[16]), .Z(n15266) );
  CND2X1 U14183 ( .A(n17787), .B(entrophy[7]), .Z(n15265) );
  CAN2X1 U14184 ( .A(n15266), .B(n15265), .Z(n15280) );
  CND2X1 U14185 ( .A(n15268), .B(n15267), .Z(n15272) );
  CND2X1 U14186 ( .A(n15348), .B(entrophy[30]), .Z(n15269) );
  CND2X1 U14187 ( .A(n15270), .B(n15269), .Z(n15271) );
  COAN1X1 U14188 ( .A(n15272), .B(n15271), .C(n12216), .Z(n15278) );
  CND3X1 U14189 ( .A(n15274), .B(datain[3]), .C(n15273), .Z(n15276) );
  CANR2XL U14190 ( .A(n17774), .B(entrophy[2]), .C(scrambler[18]), .D(n17744), 
        .Z(n15275) );
  CND2X1 U14191 ( .A(n15276), .B(n15275), .Z(n15277) );
  CNR2X1 U14192 ( .A(n15278), .B(n15277), .Z(n15279) );
  CAN3X1 U14193 ( .A(n15281), .B(n15280), .C(n15279), .Z(n15292) );
  COND1XL U14194 ( .A(n15283), .B(n15301), .C(n15282), .Z(n15285) );
  COR2X1 U14195 ( .A(n15285), .B(n15284), .Z(n15290) );
  COND1XL U14196 ( .A(n15290), .B(n15289), .C(n15288), .Z(n15291) );
  COND3X1 U14197 ( .A(n15294), .B(n15293), .C(n15292), .D(n15291), .Z(n8718)
         );
  CNR2X1 U14198 ( .A(n15296), .B(n15295), .Z(n15298) );
  COND3X1 U14199 ( .A(n15300), .B(n15299), .C(n15298), .D(n15297), .Z(n15325)
         );
  CNR2XL U14200 ( .A(n15334), .B(n15301), .Z(n15307) );
  CND3XL U14201 ( .A(n15303), .B(n15302), .C(entrophy[1]), .Z(n15304) );
  CNR2XL U14202 ( .A(n15304), .B(n17778), .Z(n15305) );
  CAOR1X1 U14203 ( .A(n15307), .B(n15306), .C(n15305), .Z(n15308) );
  CANR2XL U14204 ( .A(n15312), .B(n17804), .C(scrambler[26]), .D(n17495), .Z(
        n15316) );
  CND3X1 U14205 ( .A(n15317), .B(n15316), .C(n15315), .Z(n15324) );
  CANR1X1 U14206 ( .A(entrophy[0]), .B(n11974), .C(n15318), .Z(n15320) );
  CANR11X1 U14207 ( .A(n15322), .B(n15321), .C(n15320), .D(n12055), .Z(n15323)
         );
  CANR3X1 U14208 ( .A(n15145), .B(n15325), .C(n15324), .D(n15323), .Z(n15358)
         );
  CANR2X1 U14209 ( .A(n17775), .B(entrophy[28]), .C(entrophy[15]), .D(n11971), 
        .Z(n15326) );
  COND4CX1 U14210 ( .A(n15329), .B(n15328), .C(n15327), .D(n15326), .Z(n15342)
         );
  CND2X1 U14211 ( .A(n15330), .B(entrophy[16]), .Z(n15331) );
  COND11X1 U14212 ( .A(n15334), .B(n15333), .C(n15332), .D(n15331), .Z(n15341)
         );
  COR2XL U14213 ( .A(n15336), .B(n15335), .Z(n15337) );
  COND1XL U14214 ( .A(n15339), .B(n15338), .C(n15337), .Z(n15340) );
  CNR3X1 U14215 ( .A(n15342), .B(n15341), .C(n15340), .Z(n15357) );
  CND3XL U14216 ( .A(n15345), .B(n15344), .C(n15343), .Z(n15347) );
  COND4CX1 U14217 ( .A(entrophy[11]), .B(n15348), .C(n15347), .D(n15346), .Z(
        n15356) );
  CANR4CX1 U14218 ( .A(n15352), .B(n15351), .C(n15350), .D(n15349), .Z(n15353)
         );
  CND4X1 U14219 ( .A(n15358), .B(n15357), .C(n15356), .D(n15355), .Z(n8726) );
  CENX1 U14220 ( .A(scrambler[24]), .B(scrambler[22]), .Z(n17838) );
  CEOX1 U14221 ( .A(scrambler[29]), .B(n17838), .Z(n17842) );
  CEOX1 U14222 ( .A(scrambler[21]), .B(scrambler[20]), .Z(n17907) );
  CENX1 U14223 ( .A(n17880), .B(n17907), .Z(n17883) );
  CENX1 U14224 ( .A(scrambler[26]), .B(n17883), .Z(n17834) );
  CENX1 U14225 ( .A(scrambler[18]), .B(n17834), .Z(n15359) );
  CENX1 U14226 ( .A(n17842), .B(n15359), .Z(n15360) );
  CENX1 U14227 ( .A(polydata[6]), .B(n15360), .Z(dataout[9]) );
  CIVX2 U14228 ( .A(n18176), .Z(n17661) );
  CND2X1 U14229 ( .A(n15361), .B(poly5_shifted[65]), .Z(n15363) );
  CND2XL U14230 ( .A(n17965), .B(poly5_shifted[51]), .Z(n15362) );
  COND3X1 U14231 ( .A(n15361), .B(n17661), .C(n15363), .D(n15362), .Z(n11475)
         );
  CIVX2 U14232 ( .A(n18210), .Z(n17549) );
  CND2X1 U14233 ( .A(n17935), .B(poly5_shifted[64]), .Z(n15365) );
  CND2X1 U14234 ( .A(n17642), .B(poly5_shifted[50]), .Z(n15364) );
  COND3X1 U14235 ( .A(n15378), .B(n17549), .C(n15365), .D(n15364), .Z(n11476)
         );
  CIVXL U14236 ( .A(Poly15[50]), .Z(n15367) );
  COND1XL U14237 ( .A(poly15_shifted[50]), .B(n18210), .C(n18172), .Z(n15366)
         );
  CMXI2X1 U14238 ( .A0(n15367), .A1(n15366), .S(n16565), .Z(n9587) );
  CIVXL U14239 ( .A(Poly6[18]), .Z(n15369) );
  COND1XL U14240 ( .A(poly6_shifted[18]), .B(n18210), .C(n18172), .Z(n15368)
         );
  CMXI2X1 U14241 ( .A0(n15369), .A1(n15368), .S(n16962), .Z(n9675) );
  CENX1 U14242 ( .A(Poly2[24]), .B(Poly2[64]), .Z(n15370) );
  CENX1 U14243 ( .A(n17692), .B(n15370), .Z(n15371) );
  CNR2XL U14244 ( .A(n15371), .B(n17744), .Z(n15372) );
  CANR1XL U14245 ( .A(Poly2[36]), .B(n17306), .C(n15372), .Z(n15373) );
  COND1XL U14246 ( .A(n12005), .B(n17306), .C(n15373), .Z(n8974) );
  CEOXL U14247 ( .A(Poly12[116]), .B(Poly12[20]), .Z(n15374) );
  CANR2X1 U14248 ( .A(n12598), .B(Poly12[36]), .C(n17714), .D(n15374), .Z(
        n15375) );
  COND1XL U14249 ( .A(n12005), .B(n12598), .C(n15375), .Z(n10496) );
  CEOX1 U14250 ( .A(scrambler[25]), .B(scrambler[30]), .Z(n17871) );
  CENX1 U14251 ( .A(polydata[11]), .B(n17871), .Z(n15376) );
  CENX1 U14252 ( .A(n15376), .B(scrambler[16]), .Z(n15377) );
  CENX1 U14253 ( .A(n15377), .B(n17838), .Z(dataout[4]) );
  CIVX2 U14254 ( .A(poly5_shifted[38]), .Z(n15571) );
  CEOXL U14255 ( .A(Poly9[111]), .B(Poly9[90]), .Z(n15379) );
  CANR2X1 U14256 ( .A(n12262), .B(poly9_shifted[112]), .C(n18234), .D(n15379), 
        .Z(n15380) );
  COND1XL U14257 ( .A(n11983), .B(n12262), .C(n15380), .Z(n11204) );
  CANR2X1 U14258 ( .A(n12262), .B(Poly9[113]), .C(n17755), .D(
        poly9_shifted[113]), .Z(n15381) );
  COND1XL U14259 ( .A(n17076), .B(n12262), .C(n15381), .Z(n11192) );
  CEOXL U14260 ( .A(Poly9[91]), .B(Poly9[112]), .Z(n15382) );
  CANR2X1 U14261 ( .A(n12262), .B(poly9_shifted[113]), .C(n17449), .D(n15382), 
        .Z(n15383) );
  COND1XL U14262 ( .A(n17757), .B(n12262), .C(n15383), .Z(n11203) );
  CANR2X1 U14263 ( .A(n12262), .B(Poly9[106]), .C(n18234), .D(
        poly9_shifted[106]), .Z(n15384) );
  COND1XL U14264 ( .A(n12014), .B(n12262), .C(n15384), .Z(n11199) );
  CENX1 U14265 ( .A(Poly11[47]), .B(n15385), .Z(n15386) );
  CANR2X1 U14266 ( .A(n17683), .B(Poly11[62]), .C(n17755), .D(n15386), .Z(
        n15387) );
  COND1XL U14267 ( .A(n17004), .B(n17683), .C(n15387), .Z(n11127) );
  CENX1 U14268 ( .A(Poly11[41]), .B(n15388), .Z(n15389) );
  CANR2X1 U14269 ( .A(n17683), .B(Poly11[56]), .C(n17072), .D(n15389), .Z(
        n15390) );
  COND1XL U14270 ( .A(n16179), .B(n17683), .C(n15390), .Z(n11133) );
  CEOXL U14271 ( .A(Poly11[81]), .B(Poly11[27]), .Z(n15391) );
  CANR2X1 U14272 ( .A(n17683), .B(Poly11[42]), .C(n17449), .D(n15391), .Z(
        n15392) );
  COND1XL U14273 ( .A(n12014), .B(n17747), .C(n15392), .Z(n11147) );
  CANR2XL U14274 ( .A(n18191), .B(poly1_shifted[282]), .C(n17705), .D(
        poly1_shifted[271]), .Z(n15393) );
  COND1XL U14275 ( .A(n17196), .B(n18191), .C(n15393), .Z(n9086) );
  CANR2XL U14276 ( .A(n18191), .B(poly1_shifted[274]), .C(poly1_shifted[263]), 
        .D(n18017), .Z(n15394) );
  COND1XL U14277 ( .A(n17718), .B(n18191), .C(n15394), .Z(n9094) );
  CANR2XL U14278 ( .A(n18191), .B(poly1_shifted[275]), .C(n17998), .D(
        poly1_shifted[264]), .Z(n15395) );
  COND1XL U14279 ( .A(n17163), .B(n18191), .C(n15395), .Z(n9093) );
  CANR2XL U14280 ( .A(n17574), .B(poly7_shifted[241]), .C(n16919), .D(
        poly7_shifted[229]), .Z(n15396) );
  COND1XL U14281 ( .A(n11985), .B(n17574), .C(n15396), .Z(n9875) );
  CEOXL U14282 ( .A(Poly9[93]), .B(Poly9[114]), .Z(n15397) );
  CANR2XL U14283 ( .A(n12262), .B(poly9_shifted[115]), .C(n18017), .D(n15397), 
        .Z(n15398) );
  COND1XL U14284 ( .A(n17163), .B(n12262), .C(n15398), .Z(n11201) );
  CANR2XL U14285 ( .A(n18191), .B(poly1_shifted[294]), .C(n18234), .D(
        poly1_shifted[283]), .Z(n15399) );
  COND1XL U14286 ( .A(n17741), .B(n18191), .C(n15399), .Z(n9074) );
  CENX1 U14287 ( .A(Poly10[37]), .B(Poly10[42]), .Z(n15946) );
  CEOX1 U14288 ( .A(n15946), .B(Poly10[21]), .Z(n15400) );
  CNR2XL U14289 ( .A(n17826), .B(n15400), .Z(n15401) );
  CANR1XL U14290 ( .A(Poly10[33]), .B(n17411), .C(n15401), .Z(n15402) );
  COND1XL U14291 ( .A(n17697), .B(n17411), .C(n15402), .Z(n11070) );
  CANR2X1 U14292 ( .A(n15403), .B(Poly5[120]), .C(n17620), .D(
        poly5_shifted[120]), .Z(n15404) );
  COND1XL U14293 ( .A(n16179), .B(n15405), .C(n15404), .Z(n11406) );
  CAN2XL U14294 ( .A(n18017), .B(poly13_shifted[43]), .Z(n15406) );
  CANR1XL U14295 ( .A(poly13_shifted[57]), .B(n12900), .C(n15406), .Z(n15407)
         );
  COND1XL U14296 ( .A(n16605), .B(n12900), .C(n15407), .Z(n11017) );
  CANR2X1 U14297 ( .A(n17411), .B(Poly10[42]), .C(n17538), .D(
        poly10_shifted[42]), .Z(n15408) );
  COND1XL U14298 ( .A(n12014), .B(n17411), .C(n15408), .Z(n11061) );
  CIVXL U14299 ( .A(Poly5[0]), .Z(n15411) );
  CIVDX2 U14300 ( .A(n15613), .Z0(n17932), .Z1(n17016) );
  CNR2IX1 U14301 ( .B(Poly5[111]), .A(n15673), .Z(n15409) );
  CANR1XL U14302 ( .A(n18108), .B(n17016), .C(n15409), .Z(n15410) );
  COND1XL U14303 ( .A(n15613), .B(n15411), .C(n15410), .Z(n11526) );
  CANR2X1 U14304 ( .A(n15574), .B(n11999), .C(n17538), .D(poly5_shifted[119]), 
        .Z(n15412) );
  COND1XL U14305 ( .A(n17031), .B(n15413), .C(n15412), .Z(n11407) );
  CEOXL U14306 ( .A(Poly2[50]), .B(n17685), .Z(n15414) );
  CNR2XL U14307 ( .A(n17160), .B(n15414), .Z(n15415) );
  CANR1XL U14308 ( .A(Poly2[62]), .B(n17306), .C(n15415), .Z(n15416) );
  COND1XL U14309 ( .A(n17004), .B(n17306), .C(n15416), .Z(n8948) );
  CANR2X1 U14310 ( .A(n17016), .B(n12003), .C(n17705), .D(poly5_shifted[31]), 
        .Z(n15417) );
  COND1XL U14311 ( .A(n17016), .B(n15418), .C(n15417), .Z(n11495) );
  CANR2X1 U14312 ( .A(n12900), .B(poly13_shifted[71]), .C(n18234), .D(
        poly13_shifted[57]), .Z(n15419) );
  COND1XL U14313 ( .A(n17200), .B(n12900), .C(n15419), .Z(n11003) );
  CEOXL U14314 ( .A(n17675), .B(Poly11[20]), .Z(n15420) );
  CNR2XL U14315 ( .A(n17495), .B(n15420), .Z(n15421) );
  CANR1XL U14316 ( .A(Poly11[35]), .B(n17747), .C(n15421), .Z(n15422) );
  COND1XL U14317 ( .A(n13275), .B(n17683), .C(n15422), .Z(n11154) );
  CANR2X1 U14318 ( .A(n12932), .B(poly14_shifted[296]), .C(n17560), .D(
        poly14_shifted[280]), .Z(n15423) );
  COND1XL U14319 ( .A(n16179), .B(n12932), .C(n15423), .Z(n10125) );
  CANR2X1 U14320 ( .A(n12932), .B(poly14_shifted[275]), .C(n17714), .D(
        poly14_shifted[259]), .Z(n15424) );
  COND1XL U14321 ( .A(n13275), .B(n12932), .C(n15424), .Z(n10146) );
  CANR2X1 U14322 ( .A(n12900), .B(poly13_shifted[70]), .C(n17965), .D(
        poly13_shifted[56]), .Z(n15425) );
  COND1XL U14323 ( .A(n16179), .B(n12900), .C(n15425), .Z(n11004) );
  CANR2X1 U14324 ( .A(n12900), .B(poly13_shifted[56]), .C(n17552), .D(
        poly13_shifted[42]), .Z(n15426) );
  COND1XL U14325 ( .A(n12014), .B(n12900), .C(n15426), .Z(n11018) );
  CEOXL U14326 ( .A(n17685), .B(Poly2[35]), .Z(n15427) );
  CNR2XL U14327 ( .A(n17495), .B(n15427), .Z(n15428) );
  CANR1XL U14328 ( .A(Poly2[47]), .B(n17306), .C(n15428), .Z(n15429) );
  COND1XL U14329 ( .A(n17196), .B(n17306), .C(n15429), .Z(n8963) );
  CANR2XL U14330 ( .A(n17574), .B(Poly7[239]), .C(n17535), .D(
        poly7_shifted[239]), .Z(n15430) );
  COND1XL U14331 ( .A(n17196), .B(n17574), .C(n15430), .Z(n9865) );
  CANR2XL U14332 ( .A(n17574), .B(Poly7[241]), .C(n17998), .D(
        poly7_shifted[241]), .Z(n15431) );
  COND1XL U14333 ( .A(n17076), .B(n17574), .C(n15431), .Z(n9863) );
  CANR2XL U14334 ( .A(n17574), .B(poly7_shifted[238]), .C(n17620), .D(
        poly7_shifted[226]), .Z(n15432) );
  COND1XL U14335 ( .A(n16775), .B(n17574), .C(n15432), .Z(n9878) );
  CANR2XL U14336 ( .A(n17574), .B(poly7_shifted[243]), .C(n18234), .D(
        poly7_shifted[231]), .Z(n15433) );
  COND1XL U14337 ( .A(n17718), .B(n17574), .C(n15433), .Z(n9873) );
  CANR2XL U14338 ( .A(n17574), .B(poly7_shifted[239]), .C(n17535), .D(
        poly7_shifted[227]), .Z(n15434) );
  COND1XL U14339 ( .A(n13275), .B(n17574), .C(n15434), .Z(n9877) );
  CANR2X1 U14340 ( .A(n12012), .B(poly1_shifted[100]), .C(n17552), .D(
        poly1_shifted[89]), .Z(n15435) );
  COND1XL U14341 ( .A(n17200), .B(n12012), .C(n15435), .Z(n9268) );
  CANR2X1 U14342 ( .A(n12012), .B(poly1_shifted[89]), .C(n17453), .D(
        poly1_shifted[78]), .Z(n15436) );
  COND1XL U14343 ( .A(n17699), .B(n12012), .C(n15436), .Z(n9279) );
  CANR2X1 U14344 ( .A(n12012), .B(poly1_shifted[102]), .C(n17449), .D(
        poly1_shifted[91]), .Z(n15437) );
  COND1XL U14345 ( .A(n17741), .B(n12012), .C(n15437), .Z(n9266) );
  CANR2X1 U14346 ( .A(n12012), .B(poly1_shifted[105]), .C(n18234), .D(
        poly1_shifted[94]), .Z(n15438) );
  COND1XL U14347 ( .A(n17004), .B(n12012), .C(n15438), .Z(n9263) );
  CAN2XL U14348 ( .A(n18017), .B(poly0_shifted[163]), .Z(n15439) );
  CANR1XL U14349 ( .A(Poly0[163]), .B(n17314), .C(n15439), .Z(n15440) );
  COND1XL U14350 ( .A(n17316), .B(n13275), .C(n15440), .Z(n9414) );
  CEOXL U14351 ( .A(n17738), .B(Poly2[19]), .Z(n15441) );
  CNR2XL U14352 ( .A(n17959), .B(n15441), .Z(n15442) );
  CANR1XL U14353 ( .A(Poly2[31]), .B(n12211), .C(n15442), .Z(n15443) );
  COND1XL U14354 ( .A(n17188), .B(n12211), .C(n15443), .Z(n8979) );
  CEOXL U14355 ( .A(n15971), .B(Poly2[18]), .Z(n15444) );
  CNR2XL U14356 ( .A(n17826), .B(n15444), .Z(n15445) );
  CANR1XL U14357 ( .A(Poly2[30]), .B(n12211), .C(n15445), .Z(n15446) );
  COND1XL U14358 ( .A(n17004), .B(n12211), .C(n15446), .Z(n8980) );
  CENX1 U14359 ( .A(Poly0[108]), .B(Poly0[207]), .Z(n15447) );
  COND1XL U14360 ( .A(n15447), .B(n17495), .C(n13418), .Z(n15448) );
  CMX2XL U14361 ( .A0(n15448), .A1(poly0_shifted[144]), .S(n15880), .Z(n9451)
         );
  CANR2XL U14362 ( .A(n16425), .B(poly1_shifted[110]), .C(n18234), .D(
        poly1_shifted[99]), .Z(n15449) );
  COND1XL U14363 ( .A(n13275), .B(n16425), .C(n15449), .Z(n9258) );
  CEOXL U14364 ( .A(n17675), .B(Poly11[66]), .Z(n15450) );
  CNR2XL U14365 ( .A(n17959), .B(n15450), .Z(n15451) );
  CANR1XL U14366 ( .A(Poly11[81]), .B(n15843), .C(n15451), .Z(n15452) );
  COND1XL U14367 ( .A(n17076), .B(n15843), .C(n15452), .Z(n11108) );
  CANR2X1 U14368 ( .A(n12900), .B(poly13_shifted[68]), .C(n16702), .D(
        poly13_shifted[54]), .Z(n15453) );
  COND1XL U14369 ( .A(n17001), .B(n12900), .C(n15453), .Z(n11006) );
  CANR2X1 U14370 ( .A(n12900), .B(poly13_shifted[53]), .C(n17620), .D(
        poly13_shifted[39]), .Z(n15454) );
  COND1XL U14371 ( .A(n16939), .B(n12900), .C(n15454), .Z(n11021) );
  CANR2X1 U14372 ( .A(n12932), .B(poly14_shifted[278]), .C(n16999), .D(
        poly14_shifted[262]), .Z(n15455) );
  COND1XL U14373 ( .A(n16779), .B(n12932), .C(n15455), .Z(n10143) );
  CANR2XL U14374 ( .A(n17491), .B(poly13_shifted[501]), .C(n17620), .D(
        poly13_shifted[487]), .Z(n15456) );
  COND1XL U14375 ( .A(n17718), .B(n17491), .C(n15456), .Z(n10573) );
  CANR2XL U14376 ( .A(n12175), .B(Poly8[3]), .C(n17238), .D(Poly8[85]), .Z(
        n15457) );
  COND1XL U14377 ( .A(n13275), .B(n12175), .C(n15457), .Z(n11398) );
  CENX1 U14378 ( .A(Poly8[86]), .B(Poly8[88]), .Z(n15458) );
  CENX1 U14379 ( .A(Poly8[7]), .B(n15458), .Z(n15459) );
  CANR2X1 U14380 ( .A(n12175), .B(poly8_shifted[35]), .C(n17755), .D(n15459), 
        .Z(n15460) );
  COND1XL U14381 ( .A(n17036), .B(n12175), .C(n15460), .Z(n11380) );
  CENX1 U14382 ( .A(Poly8[8]), .B(Poly8[87]), .Z(n15461) );
  CENX1 U14383 ( .A(Poly8[89]), .B(n15461), .Z(n15462) );
  CANR2X1 U14384 ( .A(n12175), .B(poly8_shifted[36]), .C(n17998), .D(n15462), 
        .Z(n15463) );
  COND1XL U14385 ( .A(n17753), .B(n12175), .C(n15463), .Z(n11379) );
  CANR2X1 U14386 ( .A(n12175), .B(Poly8[2]), .C(n17545), .D(Poly8[84]), .Z(
        n15464) );
  COND1XL U14387 ( .A(n16775), .B(n12175), .C(n15464), .Z(n11399) );
  CANR2X1 U14388 ( .A(n12175), .B(Poly8[10]), .C(n17458), .D(Poly8[92]), .Z(
        n15465) );
  COND1XL U14389 ( .A(n12014), .B(n12175), .C(n15465), .Z(n11391) );
  CEOXL U14390 ( .A(Poly12[125]), .B(Poly12[36]), .Z(n15466) );
  CANR2X1 U14391 ( .A(n12598), .B(Poly12[52]), .C(n17705), .D(n15466), .Z(
        n15467) );
  COND1XL U14392 ( .A(n17707), .B(n12598), .C(n15467), .Z(n10480) );
  CEOXL U14393 ( .A(Poly11[78]), .B(Poly11[70]), .Z(n15468) );
  CANR2X1 U14394 ( .A(n15843), .B(Poly11[85]), .C(n16919), .D(n15468), .Z(
        n15469) );
  COND1XL U14395 ( .A(n17036), .B(n15843), .C(n15469), .Z(n11104) );
  CANR2XL U14396 ( .A(n12598), .B(Poly12[59]), .C(n18017), .D(
        poly12_shifted[59]), .Z(n15470) );
  COND1XL U14397 ( .A(n17741), .B(n12598), .C(n15470), .Z(n10473) );
  CENX1 U14398 ( .A(Poly11[44]), .B(n15471), .Z(n15472) );
  CANR2X1 U14399 ( .A(n17683), .B(Poly11[59]), .C(n17755), .D(n15472), .Z(
        n15473) );
  COND1XL U14400 ( .A(n17741), .B(n17747), .C(n15473), .Z(n11130) );
  CEOXL U14401 ( .A(Poly9[17]), .B(Poly9[106]), .Z(n15474) );
  CENX1 U14402 ( .A(Poly9[109]), .B(n15474), .Z(n15475) );
  CNR2XL U14403 ( .A(n15475), .B(n17495), .Z(n15476) );
  CANR1XL U14404 ( .A(poly9_shifted[39]), .B(n17731), .C(n15476), .Z(n15477)
         );
  COND1XL U14405 ( .A(n11978), .B(n17731), .C(n15477), .Z(n11277) );
  CIVXL U14406 ( .A(n17738), .Z(n15478) );
  CANR2X1 U14407 ( .A(n12211), .B(poly2_shifted[13]), .C(n16372), .D(n15478), 
        .Z(n15479) );
  COND1XL U14408 ( .A(n17697), .B(n12211), .C(n15479), .Z(n9009) );
  CANR2XL U14409 ( .A(n17667), .B(poly13_shifted[208]), .C(n17755), .D(
        poly13_shifted[194]), .Z(n15480) );
  COND1XL U14410 ( .A(n16775), .B(n17667), .C(n15480), .Z(n10866) );
  CIVDX1 U14411 ( .A(n16387), .Z0(n13428), .Z1(n16303) );
  CANR2X1 U14412 ( .A(n17043), .B(poly13_shifted[400]), .C(n17640), .D(
        poly13_shifted[386]), .Z(n15481) );
  COND1XL U14413 ( .A(n16303), .B(n17043), .C(n15481), .Z(n10674) );
  CANR2X1 U14414 ( .A(n17043), .B(Poly13[394]), .C(n18234), .D(
        poly13_shifted[394]), .Z(n15482) );
  COND1XL U14415 ( .A(n12014), .B(n17043), .C(n15482), .Z(n10666) );
  CIVXL U14416 ( .A(poly5_shifted[53]), .Z(n15484) );
  CANR2X1 U14417 ( .A(n12942), .B(n18138), .C(n17523), .D(poly5_shifted[39]), 
        .Z(n15483) );
  COND1XL U14418 ( .A(n17047), .B(n15484), .C(n15483), .Z(n11487) );
  CANR2XL U14419 ( .A(n12210), .B(poly1_shifted[195]), .C(poly1_shifted[184]), 
        .D(n18017), .Z(n15485) );
  COND1XL U14420 ( .A(n17721), .B(n12210), .C(n15485), .Z(n9173) );
  CANR2X1 U14421 ( .A(n12262), .B(Poly9[108]), .C(n17533), .D(
        poly9_shifted[108]), .Z(n15486) );
  COND1XL U14422 ( .A(n17087), .B(n12262), .C(n15486), .Z(n11197) );
  CEOXL U14423 ( .A(Poly11[83]), .B(Poly11[29]), .Z(n15487) );
  CANR2X1 U14424 ( .A(n17683), .B(Poly11[44]), .C(n17285), .D(n15487), .Z(
        n15488) );
  COND1XL U14425 ( .A(n17087), .B(n17747), .C(n15488), .Z(n11145) );
  CANR2X1 U14426 ( .A(n15737), .B(poly3_shifted[21]), .C(n17362), .D(Poly3[77]), .Z(n15489) );
  COND1XL U14427 ( .A(n16939), .B(n15737), .C(n15489), .Z(n8933) );
  CIVX1 U14428 ( .A(poly0_shifted[119]), .Z(n15492) );
  COND2X1 U14429 ( .A(Poly0[119]), .B(n16274), .C(n15880), .D(n11999), .Z(
        n15490) );
  COND1XL U14430 ( .A(n15492), .B(n17826), .C(n15490), .Z(n9458) );
  CANR2X1 U14431 ( .A(n11984), .B(n16274), .C(n18047), .D(poly0_shifted[101]), 
        .Z(n15491) );
  COND1XL U14432 ( .A(n15492), .B(n16276), .C(n15491), .Z(n9476) );
  CANR2X1 U14433 ( .A(n17031), .B(n18241), .C(n18047), .D(poly5_shifted[117]), 
        .Z(n15493) );
  COND1XL U14434 ( .A(n15574), .B(n15494), .C(n15493), .Z(n11409) );
  CIVXL U14435 ( .A(Poly5[122]), .Z(n17924) );
  CANR2X1 U14436 ( .A(n17031), .B(n18095), .C(n16435), .D(poly5_shifted[122]), 
        .Z(n15495) );
  COND1XL U14437 ( .A(n17031), .B(n17924), .C(n15495), .Z(n11404) );
  CANR2X1 U14438 ( .A(n12900), .B(poly13_shifted[73]), .C(n18234), .D(
        poly13_shifted[59]), .Z(n15496) );
  COND1XL U14439 ( .A(n17741), .B(n12900), .C(n15496), .Z(n11001) );
  CANR2X1 U14440 ( .A(n12175), .B(Poly8[5]), .C(n17755), .D(Poly8[87]), .Z(
        n15497) );
  COND1XL U14441 ( .A(n11995), .B(n12175), .C(n15497), .Z(n11396) );
  CENX1 U14442 ( .A(Poly8[92]), .B(Poly8[94]), .Z(n15498) );
  CENX1 U14443 ( .A(Poly8[13]), .B(n15498), .Z(n15499) );
  CANR2X1 U14444 ( .A(n12175), .B(poly8_shifted[41]), .C(n18234), .D(n15499), 
        .Z(n15500) );
  COND1XL U14445 ( .A(n17741), .B(n12175), .C(n15500), .Z(n11374) );
  CANR2X1 U14446 ( .A(n12598), .B(Poly12[56]), .C(n17655), .D(
        poly12_shifted[56]), .Z(n15501) );
  COND1XL U14447 ( .A(n16179), .B(n12598), .C(n15501), .Z(n10476) );
  CANR2X1 U14448 ( .A(n17955), .B(poly9_shifted[92]), .C(n18234), .D(
        poly9_shifted[81]), .Z(n15502) );
  COND1XL U14449 ( .A(n17076), .B(n17955), .C(n15502), .Z(n11224) );
  CANR2X1 U14450 ( .A(n17955), .B(poly9_shifted[80]), .C(n17965), .D(
        poly9_shifted[69]), .Z(n15503) );
  COND1XL U14451 ( .A(n11989), .B(n17955), .C(n15503), .Z(n11236) );
  CANR2X1 U14452 ( .A(n12900), .B(poly13_shifted[51]), .C(n17668), .D(
        poly13_shifted[37]), .Z(n15504) );
  COND1XL U14453 ( .A(n11989), .B(n12900), .C(n15504), .Z(n11023) );
  CANR2X1 U14454 ( .A(n12932), .B(poly14_shifted[277]), .C(n16435), .D(
        poly14_shifted[261]), .Z(n15505) );
  COND1XL U14455 ( .A(n11987), .B(n12932), .C(n15505), .Z(n10144) );
  CANR2X1 U14456 ( .A(n12932), .B(poly14_shifted[299]), .C(n16307), .D(
        poly14_shifted[283]), .Z(n15506) );
  COND1XL U14457 ( .A(n17741), .B(n12932), .C(n15506), .Z(n10122) );
  CIVXL U14458 ( .A(poly0_shifted[115]), .Z(n15508) );
  CANR2X1 U14459 ( .A(n14361), .B(n16274), .C(n17375), .D(poly0_shifted[97]), 
        .Z(n15507) );
  COND1XL U14460 ( .A(n15508), .B(n16276), .C(n15507), .Z(n9480) );
  CANR2X1 U14461 ( .A(n12932), .B(poly14_shifted[287]), .C(n16323), .D(
        poly14_shifted[271]), .Z(n15509) );
  COND1XL U14462 ( .A(n17196), .B(n12932), .C(n15509), .Z(n10134) );
  CIVXL U14463 ( .A(poly0_shifted[116]), .Z(n15511) );
  CANR2X1 U14464 ( .A(n13428), .B(n16274), .C(n17375), .D(poly0_shifted[98]), 
        .Z(n15510) );
  COND1XL U14465 ( .A(n15511), .B(n16276), .C(n15510), .Z(n9479) );
  CIVX1 U14466 ( .A(Poly0[108]), .Z(n15513) );
  CANR2X1 U14467 ( .A(n13028), .B(n16274), .C(n17375), .D(poly0_shifted[108]), 
        .Z(n15512) );
  COND1XL U14468 ( .A(n15513), .B(n16276), .C(n15512), .Z(n9469) );
  CIVXL U14469 ( .A(Poly0[118]), .Z(n15515) );
  CANR2X1 U14470 ( .A(n18034), .B(n16274), .C(n17375), .D(poly0_shifted[118]), 
        .Z(n15514) );
  COND1XL U14471 ( .A(n15515), .B(n16276), .C(n15514), .Z(n9459) );
  CANR2X1 U14472 ( .A(n13129), .B(Poly14[165]), .C(n16919), .D(
        poly14_shifted[165]), .Z(n15516) );
  COND1XL U14473 ( .A(n11995), .B(n13129), .C(n15516), .Z(n10240) );
  CEOXL U14474 ( .A(Poly14[294]), .B(Poly14[174]), .Z(n15517) );
  CANR2X1 U14475 ( .A(n13129), .B(poly14_shifted[206]), .C(n17634), .D(n15517), 
        .Z(n15518) );
  COND1XL U14476 ( .A(n17004), .B(n13129), .C(n15518), .Z(n10215) );
  CEOXL U14477 ( .A(Poly14[291]), .B(Poly14[171]), .Z(n15519) );
  CANR2X1 U14478 ( .A(n13129), .B(poly14_shifted[203]), .C(n17755), .D(n15519), 
        .Z(n15520) );
  COND1XL U14479 ( .A(n17741), .B(n13129), .C(n15520), .Z(n10218) );
  CANR2X1 U14480 ( .A(n13129), .B(Poly14[170]), .C(n17714), .D(
        poly14_shifted[170]), .Z(n15521) );
  COND1XL U14481 ( .A(n12014), .B(n13129), .C(n15521), .Z(n10235) );
  CEOXL U14482 ( .A(Poly12[115]), .B(Poly12[114]), .Z(n15522) );
  CENX1 U14483 ( .A(Poly12[55]), .B(n15522), .Z(n15523) );
  CNR2XL U14484 ( .A(n15523), .B(n17829), .Z(n15524) );
  CANR1XL U14485 ( .A(poly12_shifted[87]), .B(n12161), .C(n15524), .Z(n15525)
         );
  COND1XL U14486 ( .A(n16939), .B(n12161), .C(n15525), .Z(n10461) );
  CEOXL U14487 ( .A(Poly12[116]), .B(Poly12[117]), .Z(n15526) );
  CENX1 U14488 ( .A(Poly12[57]), .B(n15526), .Z(n15527) );
  CNR2XL U14489 ( .A(n15527), .B(n17744), .Z(n15528) );
  CANR1XL U14490 ( .A(poly12_shifted[89]), .B(n12161), .C(n15528), .Z(n15529)
         );
  COND1XL U14491 ( .A(n17208), .B(n12161), .C(n15529), .Z(n10459) );
  CEOXL U14492 ( .A(n15844), .B(Poly11[18]), .Z(n15530) );
  CNR2XL U14493 ( .A(n17959), .B(n15530), .Z(n15531) );
  CANR1XL U14494 ( .A(Poly11[33]), .B(n17683), .C(n15531), .Z(n15532) );
  COND1XL U14495 ( .A(n17697), .B(n17747), .C(n15532), .Z(n11156) );
  CENX1 U14496 ( .A(n17233), .B(Poly11[85]), .Z(n15859) );
  CENX1 U14497 ( .A(Poly11[55]), .B(n15859), .Z(n15533) );
  CANR2X1 U14498 ( .A(n15843), .B(Poly11[70]), .C(n17527), .D(n15533), .Z(
        n15534) );
  COND1XL U14499 ( .A(n17757), .B(n15843), .C(n15534), .Z(n11119) );
  CANR2X1 U14500 ( .A(n17610), .B(poly1_shifted[148]), .C(n17613), .D(
        poly1_shifted[137]), .Z(n15535) );
  COND1XL U14501 ( .A(n17208), .B(n17610), .C(n15535), .Z(n9220) );
  CANR2X1 U14502 ( .A(n17610), .B(poly1_shifted[160]), .C(n17280), .D(
        poly1_shifted[149]), .Z(n15536) );
  COND1XL U14503 ( .A(n12006), .B(n17610), .C(n15536), .Z(n9208) );
  CANR2X1 U14504 ( .A(n17610), .B(poly1_shifted[154]), .C(n18234), .D(
        poly1_shifted[143]), .Z(n15537) );
  COND1XL U14505 ( .A(n17196), .B(n17610), .C(n15537), .Z(n9214) );
  CANR2X1 U14506 ( .A(n17610), .B(Poly1[158]), .C(n18234), .D(
        poly1_shifted[158]), .Z(n15538) );
  COND1XL U14507 ( .A(n17004), .B(n17610), .C(n15538), .Z(n9199) );
  CEOXL U14508 ( .A(n15645), .B(dataselector[32]), .Z(n15540) );
  CANR2X1 U14509 ( .A(n18138), .B(n18248), .C(n15710), .D(dataselector[39]), 
        .Z(n15539) );
  COND1XL U14510 ( .A(n17744), .B(n15540), .C(n15539), .Z(n8756) );
  CEOXL U14511 ( .A(dataselector[58]), .B(dataselector[62]), .Z(n15541) );
  CENX1 U14512 ( .A(dataselector[26]), .B(n15541), .Z(n15543) );
  CANR2X1 U14513 ( .A(n12020), .B(n18248), .C(n15710), .D(dataselector[33]), 
        .Z(n15542) );
  COND1XL U14514 ( .A(n15543), .B(n17495), .C(n15542), .Z(n8762) );
  CANR2X1 U14515 ( .A(n12185), .B(Poly11[30]), .C(n17755), .D(
        poly11_shifted[30]), .Z(n15544) );
  COND1XL U14516 ( .A(n17004), .B(n12185), .C(n15544), .Z(n11159) );
  CANR2X1 U14517 ( .A(n12185), .B(poly11_shifted[30]), .C(n17755), .D(
        poly11_shifted[15]), .Z(n15545) );
  COND1XL U14518 ( .A(n17196), .B(n12185), .C(n15545), .Z(n11174) );
  CAN2XL U14519 ( .A(n18017), .B(Poly11[83]), .Z(n15546) );
  CANR1XL U14520 ( .A(poly11_shifted[27]), .B(n12185), .C(n15546), .Z(n15547)
         );
  COND1XL U14521 ( .A(n17087), .B(n12185), .C(n15547), .Z(n11177) );
  CANR2X1 U14522 ( .A(n12185), .B(Poly11[22]), .C(n17552), .D(
        poly11_shifted[22]), .Z(n15548) );
  COND1XL U14523 ( .A(n17753), .B(n12185), .C(n15548), .Z(n11167) );
  CIVXL U14524 ( .A(n15844), .Z(n15549) );
  CANR2X1 U14525 ( .A(n12185), .B(poly11_shifted[16]), .C(n18234), .D(n15549), 
        .Z(n15550) );
  COND1XL U14526 ( .A(n17697), .B(n12185), .C(n15550), .Z(n11188) );
  CIVXL U14527 ( .A(n17680), .Z(n15551) );
  CANR2X1 U14528 ( .A(n12185), .B(poly11_shifted[17]), .C(n18234), .D(n15551), 
        .Z(n15552) );
  COND1XL U14529 ( .A(n16303), .B(n12185), .C(n15552), .Z(n11187) );
  CANR2X1 U14530 ( .A(n12185), .B(poly11_shifted[25]), .C(n16479), .D(
        Poly11[81]), .Z(n15553) );
  COND1XL U14531 ( .A(n12014), .B(n12185), .C(n15553), .Z(n11179) );
  CANR2X1 U14532 ( .A(n12185), .B(poly11_shifted[20]), .C(n17755), .D(n17233), 
        .Z(n15554) );
  COND1XL U14533 ( .A(n11981), .B(n12185), .C(n15554), .Z(n11184) );
  CANR2X1 U14534 ( .A(n12185), .B(Poly11[17]), .C(n17398), .D(
        poly11_shifted[17]), .Z(n15555) );
  COND1XL U14535 ( .A(n17076), .B(n12185), .C(n15555), .Z(n11172) );
  CANR2X1 U14536 ( .A(n17750), .B(Poly8[78]), .C(n17642), .D(poly8_shifted[78]), .Z(n15556) );
  COND1XL U14537 ( .A(n17699), .B(n17750), .C(n15556), .Z(n11323) );
  CEOXL U14538 ( .A(Poly8[87]), .B(Poly8[72]), .Z(n15557) );
  CANR2X1 U14539 ( .A(n17750), .B(Poly8[86]), .C(n17334), .D(n15557), .Z(
        n15558) );
  COND1XL U14540 ( .A(n17753), .B(n17750), .C(n15558), .Z(n11315) );
  CANR2X1 U14541 ( .A(n17750), .B(poly8_shifted[79]), .C(n17755), .D(
        poly8_shifted[65]), .Z(n15559) );
  COND1XL U14542 ( .A(n17711), .B(n17750), .C(n15559), .Z(n11336) );
  CEOXL U14543 ( .A(Poly8[74]), .B(Poly8[89]), .Z(n15560) );
  CANR2X1 U14544 ( .A(n17750), .B(Poly8[88]), .C(n16502), .D(n15560), .Z(
        n15561) );
  COND1XL U14545 ( .A(n17721), .B(n17750), .C(n15561), .Z(n11313) );
  CANR2X1 U14546 ( .A(n17750), .B(Poly8[76]), .C(n17620), .D(poly8_shifted[76]), .Z(n15562) );
  COND1XL U14547 ( .A(n17218), .B(n17750), .C(n15562), .Z(n11325) );
  CANR2X1 U14548 ( .A(n12932), .B(poly14_shifted[289]), .C(n16427), .D(
        poly14_shifted[273]), .Z(n15563) );
  COND1XL U14549 ( .A(n17173), .B(n12932), .C(n15563), .Z(n10132) );
  CANR2X1 U14550 ( .A(n18191), .B(poly1_shifted[292]), .C(n17449), .D(
        poly1_shifted[281]), .Z(n15564) );
  COND1XL U14551 ( .A(n17123), .B(n18191), .C(n15564), .Z(n9076) );
  CEOXL U14552 ( .A(Poly14[288]), .B(Poly14[168]), .Z(n15565) );
  CANR2X1 U14553 ( .A(n13129), .B(poly14_shifted[200]), .C(n16427), .D(n15565), 
        .Z(n15566) );
  COND1XL U14554 ( .A(n17721), .B(n13129), .C(n15566), .Z(n10221) );
  CANR2XL U14555 ( .A(n17942), .B(poly5_shifted[88]), .C(n17238), .D(
        poly5_shifted[74]), .Z(n15567) );
  COND1XL U14556 ( .A(n12014), .B(n17942), .C(n15567), .Z(n11452) );
  CANR2X1 U14557 ( .A(n13129), .B(poly14_shifted[178]), .C(n16427), .D(
        poly14_shifted[162]), .Z(n15568) );
  COND1XL U14558 ( .A(n16775), .B(n13129), .C(n15568), .Z(n10243) );
  CANR2X1 U14559 ( .A(n12185), .B(Poly11[27]), .C(n17401), .D(
        poly11_shifted[27]), .Z(n15569) );
  COND1XL U14560 ( .A(n17741), .B(n12185), .C(n15569), .Z(n11162) );
  CANR2X1 U14561 ( .A(n17016), .B(n13994), .C(n17238), .D(poly5_shifted[24]), 
        .Z(n15570) );
  COND1XL U14562 ( .A(n17016), .B(n15571), .C(n15570), .Z(n11502) );
  CANR2X1 U14563 ( .A(n15574), .B(n18034), .C(n17362), .D(poly5_shifted[118]), 
        .Z(n15572) );
  COND1XL U14564 ( .A(n15574), .B(n15573), .C(n15572), .Z(n11408) );
  CAN2XL U14565 ( .A(n18017), .B(poly13_shifted[16]), .Z(n15575) );
  CANR1XL U14566 ( .A(poly13_shifted[30]), .B(n13124), .C(n15575), .Z(n15576)
         );
  COND1XL U14567 ( .A(n17062), .B(n13124), .C(n15576), .Z(n11044) );
  CNR2IXL U14568 ( .B(Poly13[515]), .A(n17160), .Z(n15577) );
  CANR1XL U14569 ( .A(poly13_shifted[15]), .B(n13124), .C(n15577), .Z(n15578)
         );
  COND1XL U14570 ( .A(n16950), .B(n13124), .C(n15578), .Z(n11059) );
  CNR2IXL U14571 ( .B(Poly13[527]), .A(n17160), .Z(n15579) );
  CANR1XL U14572 ( .A(poly13_shifted[27]), .B(n13124), .C(n15579), .Z(n15580)
         );
  COND1XL U14573 ( .A(n17065), .B(n13124), .C(n15580), .Z(n11047) );
  CAN2XL U14574 ( .A(n18017), .B(poly13_shifted[25]), .Z(n15581) );
  CANR1XL U14575 ( .A(poly13_shifted[39]), .B(n13124), .C(n15581), .Z(n15582)
         );
  COND1XL U14576 ( .A(n17200), .B(n13124), .C(n15582), .Z(n11035) );
  CANR2X1 U14577 ( .A(n17430), .B(Poly13[522]), .C(n17634), .D(
        poly13_shifted[522]), .Z(n15584) );
  COND1XL U14578 ( .A(n12014), .B(n17430), .C(n15584), .Z(n10538) );
  CANR2X1 U14579 ( .A(n17430), .B(Poly13[527]), .C(n16427), .D(
        poly13_shifted[527]), .Z(n15585) );
  COND1XL U14580 ( .A(n17196), .B(n17430), .C(n15585), .Z(n10533) );
  CANR2X1 U14581 ( .A(n17430), .B(Poly13[524]), .C(n17401), .D(
        poly13_shifted[524]), .Z(n15586) );
  COND1XL U14582 ( .A(n17087), .B(n17430), .C(n15586), .Z(n10536) );
  CANR2X1 U14583 ( .A(n17430), .B(poly13_shifted[527]), .C(n17094), .D(
        poly13_shifted[513]), .Z(n15587) );
  COND1XL U14584 ( .A(n16950), .B(n17430), .C(n15587), .Z(n10547) );
  CANR2X1 U14585 ( .A(n12008), .B(poly14_shifted[168]), .C(n16540), .D(
        poly14_shifted[152]), .Z(n15588) );
  COND1XL U14586 ( .A(n16179), .B(n12008), .C(n15588), .Z(n10253) );
  CANR2X1 U14587 ( .A(n12008), .B(poly14_shifted[146]), .C(n17527), .D(
        poly14_shifted[130]), .Z(n15589) );
  COND1XL U14588 ( .A(n16775), .B(n12008), .C(n15589), .Z(n10275) );
  CANR2X1 U14589 ( .A(n12008), .B(poly14_shifted[159]), .C(n17535), .D(
        poly14_shifted[143]), .Z(n15590) );
  COND1XL U14590 ( .A(n17196), .B(n12008), .C(n15590), .Z(n10262) );
  CANR2X1 U14591 ( .A(n12008), .B(poly14_shifted[171]), .C(n16427), .D(
        poly14_shifted[155]), .Z(n15591) );
  COND1XL U14592 ( .A(n17741), .B(n12008), .C(n15591), .Z(n10250) );
  CANR2X1 U14593 ( .A(n12008), .B(poly14_shifted[169]), .C(n16427), .D(
        poly14_shifted[153]), .Z(n15592) );
  COND1XL U14594 ( .A(n17123), .B(n12008), .C(n15592), .Z(n10252) );
  CANR2X1 U14595 ( .A(n12008), .B(poly14_shifted[147]), .C(n17620), .D(
        poly14_shifted[131]), .Z(n15593) );
  COND1XL U14596 ( .A(n13275), .B(n12008), .C(n15593), .Z(n10274) );
  CANR2X1 U14597 ( .A(n12008), .B(poly14_shifted[174]), .C(n16644), .D(
        poly14_shifted[158]), .Z(n15594) );
  COND1XL U14598 ( .A(n17004), .B(n12008), .C(n15594), .Z(n10247) );
  CANR2X1 U14599 ( .A(n12008), .B(poly14_shifted[154]), .C(n18234), .D(
        poly14_shifted[138]), .Z(n15595) );
  COND1XL U14600 ( .A(n12014), .B(n12008), .C(n15595), .Z(n10267) );
  CANR2X1 U14601 ( .A(n12008), .B(poly14_shifted[164]), .C(n17552), .D(
        poly14_shifted[148]), .Z(n15596) );
  COND1XL U14602 ( .A(n16391), .B(n12008), .C(n15596), .Z(n10257) );
  CANR2XL U14603 ( .A(n17471), .B(poly7_shifted[96]), .C(n17215), .D(
        poly7_shifted[84]), .Z(n15597) );
  COND1XL U14604 ( .A(n16391), .B(n17471), .C(n15597), .Z(n10020) );
  CIVXL U14605 ( .A(Poly0[111]), .Z(n15599) );
  CANR2X1 U14606 ( .A(n18206), .B(n16274), .C(n17375), .D(poly0_shifted[111]), 
        .Z(n15598) );
  COND1XL U14607 ( .A(n15599), .B(n16276), .C(n15598), .Z(n9466) );
  CENX1 U14608 ( .A(dataselector[60]), .B(n16384), .Z(n18238) );
  CENX1 U14609 ( .A(dataselector[40]), .B(n18238), .Z(n15601) );
  CANR2XL U14610 ( .A(n18206), .B(n18248), .C(n15710), .D(dataselector[47]), 
        .Z(n15600) );
  COND1XL U14611 ( .A(n17744), .B(n15601), .C(n15600), .Z(n8748) );
  CEOXL U14612 ( .A(dataselector[37]), .B(n18233), .Z(n15603) );
  CANR2X1 U14613 ( .A(n16350), .B(dataselector[44]), .C(n13028), .D(n18248), 
        .Z(n15602) );
  COND1XL U14614 ( .A(n17829), .B(n15603), .C(n15602), .Z(n8751) );
  CANR2X1 U14615 ( .A(n12192), .B(Poly1[231]), .C(n17755), .D(
        poly1_shifted[231]), .Z(n15604) );
  COND1XL U14616 ( .A(n17718), .B(n12192), .C(n15604), .Z(n9126) );
  CANR2X1 U14617 ( .A(n12012), .B(poly1_shifted[88]), .C(n17642), .D(
        poly1_shifted[77]), .Z(n15605) );
  COND1XL U14618 ( .A(n17090), .B(n12012), .C(n15605), .Z(n9280) );
  CANR2X1 U14619 ( .A(n12009), .B(poly14_shifted[117]), .C(n17620), .D(
        poly14_shifted[101]), .Z(n15606) );
  COND1XL U14620 ( .A(n11987), .B(n12009), .C(n15606), .Z(n10304) );
  CANR2X1 U14621 ( .A(n12009), .B(poly14_shifted[127]), .C(n17535), .D(
        poly14_shifted[111]), .Z(n15607) );
  COND1XL U14622 ( .A(n17196), .B(n12009), .C(n15607), .Z(n10294) );
  CANR2X1 U14623 ( .A(n12009), .B(poly14_shifted[114]), .C(n17527), .D(
        poly14_shifted[98]), .Z(n15608) );
  COND1XL U14624 ( .A(n16775), .B(n12009), .C(n15608), .Z(n10307) );
  CANR2X1 U14625 ( .A(n12009), .B(poly14_shifted[115]), .C(n17527), .D(
        poly14_shifted[99]), .Z(n15609) );
  COND1XL U14626 ( .A(n13275), .B(n12009), .C(n15609), .Z(n10306) );
  CANR2X1 U14627 ( .A(n12009), .B(poly14_shifted[142]), .C(n16644), .D(
        poly14_shifted[126]), .Z(n15610) );
  COND1XL U14628 ( .A(n17004), .B(n12009), .C(n15610), .Z(n10279) );
  CANR2X1 U14629 ( .A(n12009), .B(poly14_shifted[136]), .C(n16540), .D(
        poly14_shifted[120]), .Z(n15611) );
  COND1XL U14630 ( .A(n16179), .B(n12009), .C(n15611), .Z(n10285) );
  CANR2X1 U14631 ( .A(n12009), .B(poly14_shifted[139]), .C(n17063), .D(
        poly14_shifted[123]), .Z(n15612) );
  COND1XL U14632 ( .A(n17741), .B(n12009), .C(n15612), .Z(n10282) );
  CIVXL U14633 ( .A(Poly5[3]), .Z(n15615) );
  CANR2XL U14634 ( .A(n15613), .B(n18053), .C(n17714), .D(Poly5[114]), .Z(
        n15614) );
  COND1XL U14635 ( .A(n17016), .B(n15615), .C(n15614), .Z(n11523) );
  CAN2XL U14636 ( .A(n18017), .B(poly13_shifted[41]), .Z(n15616) );
  CANR1XL U14637 ( .A(poly13_shifted[55]), .B(n12900), .C(n15616), .Z(n15617)
         );
  COND1XL U14638 ( .A(n12002), .B(n12900), .C(n15617), .Z(n11019) );
  CEOXL U14639 ( .A(Poly9[94]), .B(Poly9[115]), .Z(n15618) );
  CANR2X1 U14640 ( .A(n12262), .B(Poly9[105]), .C(n17535), .D(n15618), .Z(
        n15619) );
  COND1XL U14641 ( .A(n12002), .B(n12262), .C(n15619), .Z(n11200) );
  CANR2X1 U14642 ( .A(n17731), .B(poly9_shifted[13]), .C(n17063), .D(
        Poly9[107]), .Z(n15620) );
  COND1XL U14643 ( .A(n16775), .B(n17731), .C(n15620), .Z(n11303) );
  CANR2X1 U14644 ( .A(n17731), .B(poly9_shifted[23]), .C(n17705), .D(
        poly9_shifted[12]), .Z(n15621) );
  COND1XL U14645 ( .A(n17218), .B(n17731), .C(n15621), .Z(n11293) );
  CANR2X1 U14646 ( .A(n17731), .B(Poly9[17]), .C(n17613), .D(poly9_shifted[17]), .Z(n15622) );
  COND1XL U14647 ( .A(n17076), .B(n17731), .C(n15622), .Z(n11288) );
  CANR2X1 U14648 ( .A(n17731), .B(poly9_shifted[21]), .C(n18047), .D(
        Poly9[115]), .Z(n15623) );
  COND1XL U14649 ( .A(n12014), .B(n17731), .C(n15623), .Z(n11295) );
  CEOXL U14650 ( .A(Poly9[105]), .B(Poly9[13]), .Z(n15624) );
  CANR2X1 U14651 ( .A(n17731), .B(Poly9[24]), .C(n17620), .D(n15624), .Z(
        n15625) );
  COND1XL U14652 ( .A(n16179), .B(n17731), .C(n15625), .Z(n11281) );
  CANR2X1 U14653 ( .A(n17955), .B(poly9_shifted[84]), .C(n18234), .D(
        poly9_shifted[73]), .Z(n15626) );
  COND1XL U14654 ( .A(n12002), .B(n17955), .C(n15626), .Z(n11232) );
  CANR2XL U14655 ( .A(n17491), .B(poly13_shifted[503]), .C(n17998), .D(
        poly13_shifted[489]), .Z(n15627) );
  COND1XL U14656 ( .A(n12002), .B(n17491), .C(n15627), .Z(n10571) );
  CEOXL U14657 ( .A(Poly11[80]), .B(Poly11[26]), .Z(n15628) );
  CANR2X1 U14658 ( .A(n17683), .B(Poly11[41]), .C(n16323), .D(n15628), .Z(
        n15629) );
  COND1XL U14659 ( .A(n12002), .B(n17683), .C(n15629), .Z(n11148) );
  CANR2X1 U14660 ( .A(n17731), .B(Poly9[16]), .C(n17398), .D(poly9_shifted[16]), .Z(n15630) );
  COND1XL U14661 ( .A(n17062), .B(n17731), .C(n15630), .Z(n11289) );
  CANR2XL U14662 ( .A(n16425), .B(poly1_shifted[123]), .C(n17206), .D(
        poly1_shifted[112]), .Z(n15631) );
  COND1XL U14663 ( .A(n17062), .B(n16425), .C(n15631), .Z(n9245) );
  CEOXL U14664 ( .A(Poly8[92]), .B(Poly8[77]), .Z(n15632) );
  CANR2X1 U14665 ( .A(n17750), .B(Poly8[91]), .C(n17245), .D(n15632), .Z(
        n15633) );
  COND1XL U14666 ( .A(n17741), .B(n17750), .C(n15633), .Z(n11310) );
  CANR2X1 U14667 ( .A(n17750), .B(Poly8[70]), .C(n17453), .D(poly8_shifted[70]), .Z(n15634) );
  COND1XL U14668 ( .A(n17757), .B(n17750), .C(n15634), .Z(n11331) );
  CEOXL U14669 ( .A(Poly8[95]), .B(Poly8[80]), .Z(n15635) );
  CANR2X1 U14670 ( .A(n17750), .B(Poly8[94]), .C(n18234), .D(n15635), .Z(
        n15636) );
  COND1XL U14671 ( .A(n17004), .B(n17750), .C(n15636), .Z(n11307) );
  CANR2X1 U14672 ( .A(n17750), .B(Poly8[74]), .C(n18234), .D(poly8_shifted[74]), .Z(n15637) );
  COND1XL U14673 ( .A(n12014), .B(n17750), .C(n15637), .Z(n11327) );
  CANR2X1 U14674 ( .A(n17750), .B(Poly8[69]), .C(n17348), .D(poly8_shifted[69]), .Z(n15638) );
  COND1XL U14675 ( .A(n11989), .B(n17750), .C(n15638), .Z(n11332) );
  CEOXL U14676 ( .A(n15640), .B(n15639), .Z(n15641) );
  CNR2XL U14677 ( .A(n15641), .B(n17744), .Z(n15642) );
  CANR1XL U14678 ( .A(poly4_shifted[24]), .B(n18230), .C(n15642), .Z(n15643)
         );
  COND1XL U14679 ( .A(n16939), .B(n18230), .C(n15643), .Z(n8849) );
  CENX1 U14680 ( .A(dataselector[62]), .B(dataselector[55]), .Z(n15644) );
  CENX1 U14681 ( .A(n15645), .B(n15644), .Z(n15647) );
  CANR2XL U14682 ( .A(n18105), .B(n18248), .C(n15710), .D(dataselector[62]), 
        .Z(n15646) );
  COND1XL U14683 ( .A(n15648), .B(n15647), .C(n15646), .Z(n8733) );
  CANR2X1 U14684 ( .A(n17615), .B(poly13_shifted[329]), .C(n17755), .D(
        poly13_shifted[315]), .Z(n15649) );
  COND1XL U14685 ( .A(n17741), .B(n17615), .C(n15649), .Z(n10745) );
  CEOXL U14686 ( .A(n15651), .B(n15650), .Z(n15652) );
  CNR2XL U14687 ( .A(n15652), .B(n17495), .Z(n15653) );
  CANR1XL U14688 ( .A(poly4_shifted[27]), .B(n18230), .C(n15653), .Z(n15654)
         );
  COND1XL U14689 ( .A(n12014), .B(n18230), .C(n15654), .Z(n8846) );
  CEOXL U14690 ( .A(Poly7[407]), .B(Poly7[241]), .Z(n15655) );
  CANR2XL U14691 ( .A(n17574), .B(poly7_shifted[265]), .C(n17634), .D(n15655), 
        .Z(n15656) );
  COND1XL U14692 ( .A(n17185), .B(n17574), .C(n15656), .Z(n9851) );
  CANR2X1 U14693 ( .A(n12008), .B(poly14_shifted[173]), .C(n17545), .D(
        poly14_shifted[157]), .Z(n15657) );
  COND1XL U14694 ( .A(n17185), .B(n12008), .C(n15657), .Z(n10248) );
  CANR2XL U14695 ( .A(n17667), .B(poly13_shifted[235]), .C(n16700), .D(
        poly13_shifted[221]), .Z(n15658) );
  COND1XL U14696 ( .A(n17185), .B(n17667), .C(n15658), .Z(n10839) );
  CAN2XL U14697 ( .A(n18017), .B(poly11_shifted[29]), .Z(n15659) );
  CANR1XL U14698 ( .A(Poly11[29]), .B(n12185), .C(n15659), .Z(n15660) );
  COND1XL U14699 ( .A(n17185), .B(n12185), .C(n15660), .Z(n11160) );
  CANR2X1 U14700 ( .A(n12598), .B(Poly12[61]), .C(n17755), .D(
        poly12_shifted[61]), .Z(n15661) );
  COND1XL U14701 ( .A(n17185), .B(n12598), .C(n15661), .Z(n10471) );
  CEOXL U14702 ( .A(Poly14[293]), .B(Poly14[173]), .Z(n15662) );
  CANR2X1 U14703 ( .A(n13129), .B(poly14_shifted[205]), .C(n16323), .D(n15662), 
        .Z(n15663) );
  COND1XL U14704 ( .A(n17185), .B(n13129), .C(n15663), .Z(n10216) );
  CEOXL U14705 ( .A(Poly8[94]), .B(Poly8[79]), .Z(n15664) );
  CANR2X1 U14706 ( .A(n17750), .B(Poly8[93]), .C(n18234), .D(n15664), .Z(
        n15665) );
  COND1XL U14707 ( .A(n17185), .B(n17750), .C(n15665), .Z(n11308) );
  CANR2X1 U14708 ( .A(n12900), .B(poly13_shifted[75]), .C(n16312), .D(
        poly13_shifted[61]), .Z(n15666) );
  COND1XL U14709 ( .A(n17185), .B(n12900), .C(n15666), .Z(n10999) );
  CANR2X1 U14710 ( .A(n12932), .B(Poly14[285]), .C(n17504), .D(
        poly14_shifted[285]), .Z(n15667) );
  COND1XL U14711 ( .A(n17185), .B(n12932), .C(n15667), .Z(n10120) );
  CANR2XL U14712 ( .A(n18191), .B(poly1_shifted[296]), .C(n17288), .D(
        poly1_shifted[285]), .Z(n15668) );
  COND1XL U14713 ( .A(n17185), .B(n18191), .C(n15668), .Z(n9072) );
  CANR2XL U14714 ( .A(n12009), .B(poly14_shifted[141]), .C(poly14_shifted[125]), .D(n18017), .Z(n15669) );
  COND1XL U14715 ( .A(n17185), .B(n12009), .C(n15669), .Z(n10280) );
  CANR2X1 U14716 ( .A(n12211), .B(poly2_shifted[21]), .C(n16919), .D(Poly2[67]), .Z(n15670) );
  COND1XL U14717 ( .A(n17208), .B(n12211), .C(n15670), .Z(n9001) );
  CANR2X1 U14718 ( .A(n13129), .B(Poly14[180]), .C(n17398), .D(
        poly14_shifted[180]), .Z(n15674) );
  COND1XL U14719 ( .A(n16391), .B(n13129), .C(n15674), .Z(n10225) );
  CIVX1 U14720 ( .A(Poly0[104]), .Z(n15676) );
  CANR2X1 U14721 ( .A(n18142), .B(n16274), .C(n17290), .D(poly0_shifted[104]), 
        .Z(n15675) );
  COND1XL U14722 ( .A(n15676), .B(n16276), .C(n15675), .Z(n9473) );
  CIVXL U14723 ( .A(Poly0[106]), .Z(n15678) );
  CANR2XL U14724 ( .A(n12013), .B(n16274), .C(n17290), .D(poly0_shifted[106]), 
        .Z(n15677) );
  COND1XL U14725 ( .A(n15678), .B(n16276), .C(n15677), .Z(n9471) );
  CIVXL U14726 ( .A(Poly0[107]), .Z(n15680) );
  CANR2X1 U14727 ( .A(n16381), .B(n16274), .C(n17290), .D(poly0_shifted[107]), 
        .Z(n15679) );
  COND1XL U14728 ( .A(n15680), .B(n16276), .C(n15679), .Z(n9470) );
  CIVXL U14729 ( .A(poly0_shifted[114]), .Z(n15682) );
  CANR2X1 U14730 ( .A(n18108), .B(n16274), .C(n17290), .D(poly0_shifted[96]), 
        .Z(n15681) );
  COND1XL U14731 ( .A(n15682), .B(n16276), .C(n15681), .Z(n9481) );
  CANR2X1 U14732 ( .A(n12932), .B(poly14_shifted[300]), .C(n16919), .D(
        poly14_shifted[284]), .Z(n15683) );
  COND1XL U14733 ( .A(n11978), .B(n12932), .C(n15683), .Z(n10121) );
  CANR2X1 U14734 ( .A(n12161), .B(Poly12[66]), .C(n17755), .D(
        poly12_shifted[66]), .Z(n15684) );
  COND1XL U14735 ( .A(n16303), .B(n12161), .C(n15684), .Z(n10466) );
  CANR2X1 U14736 ( .A(n12161), .B(Poly12[89]), .C(n17998), .D(
        poly12_shifted[89]), .Z(n15685) );
  COND1XL U14737 ( .A(n17123), .B(n12161), .C(n15685), .Z(n10443) );
  CANR2X1 U14738 ( .A(n12161), .B(Poly12[84]), .C(n17755), .D(
        poly12_shifted[84]), .Z(n15686) );
  COND1XL U14739 ( .A(n17707), .B(n12161), .C(n15686), .Z(n10448) );
  CANR2X1 U14740 ( .A(n17955), .B(poly9_shifted[85]), .C(n17538), .D(
        poly9_shifted[74]), .Z(n15687) );
  COND1XL U14741 ( .A(n12014), .B(n17955), .C(n15687), .Z(n11231) );
  CANR2XL U14742 ( .A(n17955), .B(Poly9[85]), .C(n18017), .D(poly9_shifted[85]), .Z(n15688) );
  COND1XL U14743 ( .A(n17036), .B(n17955), .C(n15688), .Z(n11220) );
  CANR2X1 U14744 ( .A(n17955), .B(Poly9[93]), .C(n17640), .D(poly9_shifted[93]), .Z(n15689) );
  COND1XL U14745 ( .A(n17185), .B(n17955), .C(n15689), .Z(n11212) );
  CIVDX1 U14746 ( .A(n17753), .Z0(n14487), .Z1(n17001) );
  CANR2X1 U14747 ( .A(n12932), .B(poly14_shifted[294]), .C(n16999), .D(
        poly14_shifted[278]), .Z(n15690) );
  COND1XL U14748 ( .A(n17001), .B(n12932), .C(n15690), .Z(n10127) );
  CAN2XL U14749 ( .A(n18017), .B(poly12_shifted[54]), .Z(n15691) );
  CANR1XL U14750 ( .A(Poly12[54]), .B(n12598), .C(n15691), .Z(n15692) );
  COND1XL U14751 ( .A(n17001), .B(n12598), .C(n15692), .Z(n10478) );
  CANR2X1 U14752 ( .A(n12009), .B(poly14_shifted[128]), .C(n17755), .D(
        poly14_shifted[112]), .Z(n15693) );
  COND1XL U14753 ( .A(n17211), .B(n12009), .C(n15693), .Z(n10293) );
  CANR2X1 U14754 ( .A(n17750), .B(Poly8[80]), .C(n17965), .D(poly8_shifted[80]), .Z(n15694) );
  COND1XL U14755 ( .A(n17211), .B(n17750), .C(n15694), .Z(n11321) );
  CANR2X1 U14756 ( .A(n12008), .B(poly14_shifted[160]), .C(n17705), .D(
        poly14_shifted[144]), .Z(n15695) );
  COND1XL U14757 ( .A(n17211), .B(n12008), .C(n15695), .Z(n10261) );
  CANR2X1 U14758 ( .A(n13129), .B(Poly14[175]), .C(n16999), .D(
        poly14_shifted[175]), .Z(n15696) );
  COND1XL U14759 ( .A(n17196), .B(n13129), .C(n15696), .Z(n10230) );
  CANR2X1 U14760 ( .A(n17615), .B(poly13_shifted[318]), .C(n17504), .D(
        poly13_shifted[304]), .Z(n15697) );
  COND1XL U14761 ( .A(n17062), .B(n17615), .C(n15697), .Z(n10756) );
  CANR2X1 U14762 ( .A(n18018), .B(poly7_shifted[24]), .C(n17105), .D(
        poly7_shifted[12]), .Z(n15698) );
  COND1XL U14763 ( .A(n17218), .B(n18018), .C(n15698), .Z(n10092) );
  CANR2X1 U14764 ( .A(n18018), .B(Poly7[21]), .C(n17535), .D(poly7_shifted[21]), .Z(n15699) );
  COND1XL U14765 ( .A(n12006), .B(n18018), .C(n15699), .Z(n10083) );
  CANR2X1 U14766 ( .A(n18018), .B(Poly7[30]), .C(n16372), .D(poly7_shifted[30]), .Z(n15700) );
  COND1XL U14767 ( .A(n17004), .B(n17564), .C(n15700), .Z(n10074) );
  CANR2X1 U14768 ( .A(n13124), .B(poly13_shifted[28]), .C(n17705), .D(
        poly13_shifted[14]), .Z(n15701) );
  COND1XL U14769 ( .A(n17699), .B(n13124), .C(n15701), .Z(n11046) );
  CANR2X1 U14770 ( .A(n13124), .B(poly13_shifted[34]), .C(n17504), .D(
        poly13_shifted[20]), .Z(n15702) );
  COND1XL U14771 ( .A(n17707), .B(n13124), .C(n15702), .Z(n11040) );
  CANR2X1 U14772 ( .A(n13124), .B(poly13_shifted[41]), .C(n17705), .D(
        poly13_shifted[27]), .Z(n15703) );
  COND1XL U14773 ( .A(n17741), .B(n13124), .C(n15703), .Z(n11033) );
  CIVDX1 U14774 ( .A(n16387), .Z0(n12415), .Z1(n16775) );
  CANR2X1 U14775 ( .A(n13124), .B(poly13_shifted[16]), .C(n17072), .D(
        Poly13[516]), .Z(n15704) );
  COND1XL U14776 ( .A(n16775), .B(n13124), .C(n15704), .Z(n11058) );
  CANR2X1 U14777 ( .A(n13124), .B(poly13_shifted[29]), .C(n17401), .D(
        poly13_shifted[15]), .Z(n15705) );
  COND1XL U14778 ( .A(n17196), .B(n13124), .C(n15705), .Z(n11045) );
  CANR2X1 U14779 ( .A(n13124), .B(poly13_shifted[44]), .C(n17998), .D(
        poly13_shifted[30]), .Z(n15706) );
  COND1XL U14780 ( .A(n13418), .B(n13124), .C(n15706), .Z(n11030) );
  CANR2XL U14781 ( .A(n13124), .B(poly13_shifted[26]), .C(n17998), .D(
        Poly13[526]), .Z(n15707) );
  COND1XL U14782 ( .A(n17087), .B(n13124), .C(n15707), .Z(n11048) );
  CANR2X1 U14783 ( .A(n13124), .B(poly13_shifted[36]), .C(n17755), .D(
        poly13_shifted[22]), .Z(n15708) );
  COND1XL U14784 ( .A(n17001), .B(n13124), .C(n15708), .Z(n11038) );
  CEOXL U14785 ( .A(dataselector[33]), .B(n17821), .Z(n15709) );
  CENX1 U14786 ( .A(n15981), .B(n15709), .Z(n15712) );
  CANR2X1 U14787 ( .A(n18142), .B(n18248), .C(n15710), .D(dataselector[40]), 
        .Z(n15711) );
  COND1XL U14788 ( .A(n17495), .B(n15712), .C(n15711), .Z(n8755) );
  CEOXL U14789 ( .A(Poly7[399]), .B(Poly7[233]), .Z(n15713) );
  CANR2X1 U14790 ( .A(n17574), .B(poly7_shifted[257]), .C(n16985), .D(n15713), 
        .Z(n15714) );
  COND1XL U14791 ( .A(n12006), .B(n17574), .C(n15714), .Z(n9859) );
  CANR2X1 U14792 ( .A(n17574), .B(Poly7[237]), .C(n16488), .D(
        poly7_shifted[237]), .Z(n15715) );
  COND1XL U14793 ( .A(n17090), .B(n17574), .C(n15715), .Z(n9867) );
  CEOXL U14794 ( .A(Poly7[405]), .B(Poly7[239]), .Z(n15716) );
  CANR2X1 U14795 ( .A(n17574), .B(poly7_shifted[263]), .C(n17401), .D(n15716), 
        .Z(n15717) );
  COND1XL U14796 ( .A(n17741), .B(n17574), .C(n15717), .Z(n9853) );
  CANR2X1 U14797 ( .A(n17574), .B(Poly7[240]), .C(n17535), .D(
        poly7_shifted[240]), .Z(n15718) );
  COND1XL U14798 ( .A(n17211), .B(n17574), .C(n15718), .Z(n9864) );
  CANR2X1 U14799 ( .A(n12008), .B(poly14_shifted[153]), .C(n16695), .D(
        poly14_shifted[137]), .Z(n15719) );
  COND1XL U14800 ( .A(n17208), .B(n12008), .C(n15719), .Z(n10268) );
  CANR2X1 U14801 ( .A(n17430), .B(Poly13[521]), .C(n17072), .D(
        poly13_shifted[521]), .Z(n15720) );
  COND1XL U14802 ( .A(n17208), .B(n17430), .C(n15720), .Z(n10539) );
  CANR2X1 U14803 ( .A(n12932), .B(poly14_shifted[281]), .C(n17063), .D(
        poly14_shifted[265]), .Z(n15721) );
  COND1XL U14804 ( .A(n17208), .B(n12932), .C(n15721), .Z(n10140) );
  CANR2X1 U14805 ( .A(n18018), .B(poly7_shifted[21]), .C(n17535), .D(
        Poly7[408]), .Z(n15722) );
  COND1XL U14806 ( .A(n17208), .B(n18018), .C(n15722), .Z(n10095) );
  CEOXL U14807 ( .A(Poly12[114]), .B(Poly12[121]), .Z(n15723) );
  CENX1 U14808 ( .A(Poly12[25]), .B(n15723), .Z(n15724) );
  CNR2XL U14809 ( .A(n15724), .B(n17744), .Z(n15725) );
  CANR1XL U14810 ( .A(poly12_shifted[57]), .B(n12598), .C(n15725), .Z(n15726)
         );
  COND1XL U14811 ( .A(n17208), .B(n12598), .C(n15726), .Z(n10491) );
  CANR2X1 U14812 ( .A(n17574), .B(Poly7[233]), .C(n17178), .D(
        poly7_shifted[233]), .Z(n15727) );
  COND1XL U14813 ( .A(n17208), .B(n17574), .C(n15727), .Z(n9871) );
  CANR2X1 U14814 ( .A(n12958), .B(poly14_shifted[97]), .C(n17362), .D(
        poly14_shifted[81]), .Z(n15728) );
  COND1XL U14815 ( .A(n17173), .B(n12958), .C(n15728), .Z(n10324) );
  CANR2X1 U14816 ( .A(n12958), .B(poly14_shifted[109]), .C(n17466), .D(
        poly14_shifted[93]), .Z(n15729) );
  COND1XL U14817 ( .A(n17185), .B(n12958), .C(n15729), .Z(n10312) );
  CANR2X1 U14818 ( .A(n12958), .B(poly14_shifted[83]), .C(n18234), .D(
        poly14_shifted[67]), .Z(n15730) );
  COND1XL U14819 ( .A(n13275), .B(n12958), .C(n15730), .Z(n10338) );
  CANR2X1 U14820 ( .A(n12958), .B(poly14_shifted[85]), .C(n17620), .D(
        poly14_shifted[69]), .Z(n15731) );
  COND1XL U14821 ( .A(n11981), .B(n12958), .C(n15731), .Z(n10336) );
  CANR2X1 U14822 ( .A(n12958), .B(poly14_shifted[107]), .C(n17063), .D(
        poly14_shifted[91]), .Z(n15732) );
  COND1XL U14823 ( .A(n17741), .B(n12958), .C(n15732), .Z(n10314) );
  CANR2X1 U14824 ( .A(n12958), .B(poly14_shifted[96]), .C(n17375), .D(
        poly14_shifted[80]), .Z(n15733) );
  COND1XL U14825 ( .A(n17062), .B(n12958), .C(n15733), .Z(n10325) );
  CANR2XL U14826 ( .A(n18191), .B(poly1_shifted[269]), .C(n16326), .D(
        poly1_shifted[258]), .Z(n15734) );
  COND1XL U14827 ( .A(n16775), .B(n18191), .C(n15734), .Z(n9099) );
  CANR2X1 U14828 ( .A(n18191), .B(poly1_shifted[291]), .C(n16326), .D(
        poly1_shifted[280]), .Z(n15735) );
  COND1XL U14829 ( .A(n17721), .B(n18191), .C(n15735), .Z(n9077) );
  CND2X1 U14830 ( .A(n15737), .B(poly3_shifted[26]), .Z(n15736) );
  COND4CXL U14831 ( .A(n17218), .B(n16728), .C(n15737), .D(n15736), .Z(n8928)
         );
  CANR2X1 U14832 ( .A(n17615), .B(poly13_shifted[317]), .C(poly13_shifted[303]), .D(n16947), .Z(n15738) );
  COND1XL U14833 ( .A(n17196), .B(n17615), .C(n15738), .Z(n10757) );
  CANR2X1 U14834 ( .A(n17615), .B(poly13_shifted[324]), .C(n18017), .D(
        poly13_shifted[310]), .Z(n15739) );
  COND1XL U14835 ( .A(n17001), .B(n17615), .C(n15739), .Z(n10750) );
  CANR2X1 U14836 ( .A(n17615), .B(poly13_shifted[332]), .C(n17965), .D(
        poly13_shifted[318]), .Z(n15740) );
  COND1XL U14837 ( .A(n13418), .B(n17615), .C(n15740), .Z(n10742) );
  CANR2X1 U14838 ( .A(n18002), .B(poly14_shifted[26]), .C(n18234), .D(
        Poly14[295]), .Z(n15741) );
  COND1XL U14839 ( .A(n12014), .B(n18002), .C(n15741), .Z(n10395) );
  CANR2X1 U14840 ( .A(n18002), .B(poly14_shifted[22]), .C(n17714), .D(
        Poly14[291]), .Z(n15742) );
  COND1XL U14841 ( .A(n16779), .B(n18002), .C(n15742), .Z(n10399) );
  CANR2X1 U14842 ( .A(n18002), .B(poly14_shifted[44]), .C(n17401), .D(
        poly14_shifted[28]), .Z(n15743) );
  COND1XL U14843 ( .A(n11978), .B(n18002), .C(n15743), .Z(n10377) );
  CANR2XL U14844 ( .A(n17332), .B(Poly1[345]), .C(n17285), .D(
        poly1_shifted[345]), .Z(n15744) );
  COND1XL U14845 ( .A(n17123), .B(n17332), .C(n15744), .Z(n9012) );
  CANR2XL U14846 ( .A(n17332), .B(Poly1[342]), .C(n17998), .D(
        poly1_shifted[342]), .Z(n15745) );
  COND1XL U14847 ( .A(n17753), .B(n17332), .C(n15745), .Z(n9015) );
  CANR2XL U14848 ( .A(n17332), .B(Poly1[344]), .C(n16326), .D(
        poly1_shifted[344]), .Z(n15746) );
  COND1XL U14849 ( .A(n17721), .B(n17332), .C(n15746), .Z(n9013) );
  CANR2X1 U14850 ( .A(n17750), .B(Poly8[77]), .C(n17174), .D(poly8_shifted[77]), .Z(n15747) );
  COND1XL U14851 ( .A(n17065), .B(n17750), .C(n15747), .Z(n11324) );
  CAN2XL U14852 ( .A(n18017), .B(poly9_shifted[109]), .Z(n15748) );
  CANR1XL U14853 ( .A(Poly9[109]), .B(n12262), .C(n15748), .Z(n15749) );
  COND1XL U14854 ( .A(n17065), .B(n12262), .C(n15749), .Z(n11196) );
  CANR2X1 U14855 ( .A(n12175), .B(Poly8[13]), .C(n17552), .D(Poly8[95]), .Z(
        n15750) );
  COND1XL U14856 ( .A(n17065), .B(n12175), .C(n15750), .Z(n11388) );
  CANR2XL U14857 ( .A(n12185), .B(poly11_shifted[28]), .C(n17705), .D(
        Poly11[84]), .Z(n15751) );
  COND1XL U14858 ( .A(n17065), .B(n12185), .C(n15751), .Z(n11176) );
  CAN2XL U14859 ( .A(n18017), .B(poly12_shifted[93]), .Z(n15752) );
  CANR1XL U14860 ( .A(Poly12[93]), .B(n12161), .C(n15752), .Z(n15753) );
  COND1XL U14861 ( .A(n17185), .B(n12161), .C(n15753), .Z(n10439) );
  CENX1 U14862 ( .A(dataselector[30]), .B(n18238), .Z(n15755) );
  CANR2X1 U14863 ( .A(n11986), .B(n18248), .C(dataselector[37]), .D(n16350), 
        .Z(n15754) );
  COND1XL U14864 ( .A(n17744), .B(n15755), .C(n15754), .Z(n8758) );
  CEOXL U14865 ( .A(Poly1[346]), .B(Poly1[208]), .Z(n15756) );
  CANR2X1 U14866 ( .A(n17053), .B(poly1_shifted[230]), .C(n17538), .D(n15756), 
        .Z(n15757) );
  COND1XL U14867 ( .A(n17741), .B(n17053), .C(n15757), .Z(n9138) );
  CANR2X1 U14868 ( .A(n17053), .B(Poly1[208]), .C(n17072), .D(
        poly1_shifted[208]), .Z(n15758) );
  COND1XL U14869 ( .A(n17062), .B(n17053), .C(n15758), .Z(n9149) );
  CANR2X1 U14870 ( .A(n17053), .B(Poly1[205]), .C(n17538), .D(
        poly1_shifted[205]), .Z(n15759) );
  COND1XL U14871 ( .A(n17090), .B(n17053), .C(n15759), .Z(n9152) );
  CANR2X1 U14872 ( .A(n17053), .B(poly1_shifted[205]), .C(n17144), .D(
        poly1_shifted[194]), .Z(n15760) );
  COND1XL U14873 ( .A(n16775), .B(n17053), .C(n15760), .Z(n9163) );
  CANR2X1 U14874 ( .A(n17053), .B(Poly1[207]), .C(n17156), .D(
        poly1_shifted[207]), .Z(n15761) );
  COND1XL U14875 ( .A(n17196), .B(n17053), .C(n15761), .Z(n9150) );
  CANR2X1 U14876 ( .A(n17731), .B(Poly9[22]), .C(n16919), .D(poly9_shifted[22]), .Z(n15762) );
  COND1XL U14877 ( .A(n17753), .B(n17731), .C(n15762), .Z(n11283) );
  CANR2X1 U14878 ( .A(n17731), .B(Poly9[15]), .C(n17620), .D(poly9_shifted[15]), .Z(n15763) );
  COND1XL U14879 ( .A(n17196), .B(n17731), .C(n15763), .Z(n11290) );
  CANR2X1 U14880 ( .A(n17731), .B(poly9_shifted[17]), .C(n16326), .D(
        Poly9[111]), .Z(n15764) );
  COND1XL U14881 ( .A(n17757), .B(n17731), .C(n15764), .Z(n11299) );
  CENX1 U14882 ( .A(Poly9[105]), .B(Poly9[108]), .Z(n15765) );
  CENX1 U14883 ( .A(Poly9[16]), .B(n15765), .Z(n15766) );
  CANR2X1 U14884 ( .A(n17731), .B(poly9_shifted[38]), .C(n17755), .D(n15766), 
        .Z(n15767) );
  COND1XL U14885 ( .A(n17741), .B(n17731), .C(n15767), .Z(n11278) );
  CENX1 U14886 ( .A(Poly9[107]), .B(Poly9[110]), .Z(n15768) );
  CENX1 U14887 ( .A(Poly9[18]), .B(n15768), .Z(n15769) );
  CANR2X1 U14888 ( .A(n17731), .B(poly9_shifted[40]), .C(n17094), .D(n15769), 
        .Z(n15770) );
  COND1XL U14889 ( .A(n17185), .B(n17731), .C(n15770), .Z(n11276) );
  CENX1 U14890 ( .A(Poly9[108]), .B(Poly9[111]), .Z(n15771) );
  CENX1 U14891 ( .A(Poly9[19]), .B(n15771), .Z(n15772) );
  CANR2X1 U14892 ( .A(n17731), .B(poly9_shifted[41]), .C(n17063), .D(n15772), 
        .Z(n15773) );
  COND1XL U14893 ( .A(n13418), .B(n17731), .C(n15773), .Z(n11275) );
  CANR2X1 U14894 ( .A(n12009), .B(poly14_shifted[125]), .C(n18234), .D(
        poly14_shifted[109]), .Z(n15774) );
  COND1XL U14895 ( .A(n17090), .B(n12009), .C(n15774), .Z(n10296) );
  CANR2X1 U14896 ( .A(n12008), .B(poly14_shifted[157]), .C(n17705), .D(
        poly14_shifted[141]), .Z(n15776) );
  COND1XL U14897 ( .A(n17065), .B(n12008), .C(n15776), .Z(n10264) );
  CANR2X1 U14898 ( .A(n17430), .B(Poly13[525]), .C(n18234), .D(
        poly13_shifted[525]), .Z(n15777) );
  COND1XL U14899 ( .A(n17065), .B(n17430), .C(n15777), .Z(n10535) );
  CANR2X1 U14900 ( .A(n12210), .B(poly1_shifted[184]), .C(n17094), .D(
        poly1_shifted[173]), .Z(n15778) );
  COND1XL U14901 ( .A(n17090), .B(n12210), .C(n15778), .Z(n9184) );
  CANR2X1 U14902 ( .A(n13129), .B(Poly14[173]), .C(n17533), .D(
        poly14_shifted[173]), .Z(n15779) );
  COND1XL U14903 ( .A(n17065), .B(n13129), .C(n15779), .Z(n10232) );
  CANR2X1 U14904 ( .A(n12211), .B(poly2_shifted[25]), .C(n17174), .D(
        poly2_shifted[13]), .Z(n15780) );
  COND1XL U14905 ( .A(n17065), .B(n12211), .C(n15780), .Z(n8997) );
  CANR2X1 U14906 ( .A(n17615), .B(poly13_shifted[315]), .C(n17298), .D(
        poly13_shifted[301]), .Z(n15781) );
  COND1XL U14907 ( .A(n17090), .B(n17615), .C(n15781), .Z(n10759) );
  CANR2X1 U14908 ( .A(n12900), .B(poly13_shifted[59]), .C(n17620), .D(
        poly13_shifted[45]), .Z(n15782) );
  COND1XL U14909 ( .A(n17090), .B(n12900), .C(n15782), .Z(n11015) );
  CEOXL U14910 ( .A(Poly11[84]), .B(Poly11[30]), .Z(n15783) );
  CANR2X1 U14911 ( .A(n17683), .B(Poly11[45]), .C(n17634), .D(n15783), .Z(
        n15784) );
  COND1XL U14912 ( .A(n17090), .B(n17683), .C(n15784), .Z(n11144) );
  CEOXL U14913 ( .A(Poly11[83]), .B(Poly11[62]), .Z(n15785) );
  CANR2X1 U14914 ( .A(n15843), .B(Poly11[77]), .C(n17449), .D(n15785), .Z(
        n15786) );
  COND1XL U14915 ( .A(n17065), .B(n15843), .C(n15786), .Z(n11112) );
  CENX1 U14916 ( .A(polydata[14]), .B(scrambler[28]), .Z(n15787) );
  CEOX1 U14917 ( .A(scrambler[25]), .B(n15787), .Z(n15789) );
  CEOX1 U14918 ( .A(scrambler[30]), .B(scrambler[20]), .Z(n17875) );
  CENX1 U14919 ( .A(n17838), .B(n17884), .Z(n17921) );
  CENX1 U14920 ( .A(scrambler[26]), .B(scrambler[16]), .Z(n17912) );
  CENX1 U14921 ( .A(n17921), .B(n17912), .Z(n17889) );
  CEOX1 U14922 ( .A(n17875), .B(n17889), .Z(n15788) );
  CENX1 U14923 ( .A(n15789), .B(n15788), .Z(dataout[1]) );
  CANR2X1 U14924 ( .A(n17592), .B(poly13_shifted[275]), .C(n17755), .D(
        poly13_shifted[261]), .Z(n15790) );
  COND1XL U14925 ( .A(n11991), .B(n17592), .C(n15790), .Z(n10799) );
  CANR2X1 U14926 ( .A(n17592), .B(poly13_shifted[277]), .C(n16700), .D(
        poly13_shifted[263]), .Z(n15791) );
  COND1XL U14927 ( .A(n17718), .B(n17592), .C(n15791), .Z(n10797) );
  CANR2X1 U14928 ( .A(n17592), .B(poly13_shifted[279]), .C(n17178), .D(
        poly13_shifted[265]), .Z(n15792) );
  COND1XL U14929 ( .A(n12002), .B(n17592), .C(n15792), .Z(n10795) );
  CANR2X1 U14930 ( .A(n17592), .B(poly13_shifted[273]), .C(n17298), .D(
        poly13_shifted[259]), .Z(n15793) );
  COND1XL U14931 ( .A(n13275), .B(n17592), .C(n15793), .Z(n10801) );
  CANR2X1 U14932 ( .A(n17592), .B(poly13_shifted[282]), .C(n17453), .D(
        poly13_shifted[268]), .Z(n15794) );
  COND1XL U14933 ( .A(n17087), .B(n17592), .C(n15794), .Z(n10792) );
  CANR2X1 U14934 ( .A(n17592), .B(Poly13[276]), .C(n17634), .D(
        poly13_shifted[276]), .Z(n15795) );
  COND1XL U14935 ( .A(n17707), .B(n17592), .C(n15795), .Z(n10784) );
  CEOX1 U14936 ( .A(dataselector[18]), .B(n16135), .Z(n15796) );
  CANR2X1 U14937 ( .A(n18249), .B(n17832), .C(n16695), .D(n15796), .Z(n15797)
         );
  COND1XL U14938 ( .A(n15799), .B(n15798), .C(n15797), .Z(n8770) );
  CANR2X1 U14939 ( .A(n18018), .B(Poly7[22]), .C(n17099), .D(poly7_shifted[22]), .Z(n15800) );
  COND1XL U14940 ( .A(n17001), .B(n18018), .C(n15800), .Z(n10082) );
  CANR2X1 U14941 ( .A(n12008), .B(poly14_shifted[165]), .C(n17620), .D(
        poly14_shifted[149]), .Z(n15801) );
  COND1XL U14942 ( .A(n12006), .B(n12008), .C(n15801), .Z(n10256) );
  CEOXL U14943 ( .A(Poly3[75]), .B(Poly3[83]), .Z(n15802) );
  CENX1 U14944 ( .A(Poly3[50]), .B(n15802), .Z(n15805) );
  CND2XL U14945 ( .A(n18108), .B(n18209), .Z(n15804) );
  CND2XL U14946 ( .A(poly3_shifted[78]), .B(n17359), .Z(n15803) );
  COND3XL U14947 ( .A(n15805), .B(n17744), .C(n15804), .D(n15803), .Z(n8876)
         );
  CANR2X1 U14948 ( .A(n17430), .B(Poly13[514]), .C(n17203), .D(
        poly13_shifted[514]), .Z(n15806) );
  COND1XL U14949 ( .A(n16775), .B(n17430), .C(n15806), .Z(n10546) );
  CANR2XL U14950 ( .A(n18191), .B(poly1_shifted[273]), .C(n17215), .D(
        poly1_shifted[262]), .Z(n15807) );
  COND1XL U14951 ( .A(n17757), .B(n18191), .C(n15807), .Z(n9095) );
  CANR2XL U14952 ( .A(n18191), .B(poly1_shifted[272]), .C(n17238), .D(
        poly1_shifted[261]), .Z(n15808) );
  COND1XL U14953 ( .A(n11991), .B(n18191), .C(n15808), .Z(n9096) );
  CANR2XL U14954 ( .A(n12932), .B(Poly14[286]), .C(n17285), .D(
        poly14_shifted[286]), .Z(n15809) );
  COND1XL U14955 ( .A(n13418), .B(n12932), .C(n15809), .Z(n10119) );
  CANR2XL U14956 ( .A(n18191), .B(poly1_shifted[284]), .C(n17288), .D(
        poly1_shifted[273]), .Z(n15810) );
  COND1XL U14957 ( .A(n17173), .B(n18191), .C(n15810), .Z(n9084) );
  CANR2X1 U14958 ( .A(n17955), .B(Poly9[91]), .C(n16985), .D(poly9_shifted[91]), .Z(n15811) );
  COND1XL U14959 ( .A(n17741), .B(n17955), .C(n15811), .Z(n11214) );
  CANR2X1 U14960 ( .A(n12012), .B(poly1_shifted[99]), .C(n17209), .D(
        poly1_shifted[88]), .Z(n15812) );
  COND1XL U14961 ( .A(n17721), .B(n12012), .C(n15812), .Z(n9269) );
  CANR2XL U14962 ( .A(n18191), .B(poly1_shifted[297]), .C(n17136), .D(
        poly1_shifted[286]), .Z(n15813) );
  COND1XL U14963 ( .A(n17004), .B(n18191), .C(n15813), .Z(n9071) );
  CANR2X1 U14964 ( .A(n17053), .B(poly1_shifted[204]), .C(n16307), .D(
        poly1_shifted[193]), .Z(n15814) );
  COND1XL U14965 ( .A(n17697), .B(n17053), .C(n15814), .Z(n9164) );
  CANR2X1 U14966 ( .A(n17053), .B(poly1_shifted[208]), .C(n18047), .D(
        poly1_shifted[197]), .Z(n15815) );
  COND1XL U14967 ( .A(n11989), .B(n17053), .C(n15815), .Z(n9160) );
  CANR2X1 U14968 ( .A(n18002), .B(poly14_shifted[33]), .C(n17121), .D(
        poly14_shifted[17]), .Z(n15816) );
  COND1XL U14969 ( .A(n17173), .B(n18002), .C(n15816), .Z(n10388) );
  CANR2X1 U14970 ( .A(n12598), .B(Poly12[60]), .C(n17449), .D(
        poly12_shifted[60]), .Z(n15817) );
  COND1XL U14971 ( .A(n11978), .B(n12598), .C(n15817), .Z(n10472) );
  CANR2X1 U14972 ( .A(n17731), .B(Poly9[13]), .C(n17545), .D(poly9_shifted[13]), .Z(n15818) );
  COND1XL U14973 ( .A(n17090), .B(n17731), .C(n15818), .Z(n11292) );
  CAN2XL U14974 ( .A(n18017), .B(poly13_shifted[28]), .Z(n15819) );
  CANR1XL U14975 ( .A(poly13_shifted[42]), .B(n13124), .C(n15819), .Z(n15820)
         );
  COND1XL U14976 ( .A(n11978), .B(n13124), .C(n15820), .Z(n11032) );
  CANR2X1 U14977 ( .A(n12211), .B(poly2_shifted[22]), .C(n17203), .D(Poly2[68]), .Z(n15821) );
  COND1XL U14978 ( .A(n12014), .B(n12211), .C(n15821), .Z(n9000) );
  CIVX1 U14979 ( .A(n15822), .Z(n15823) );
  CANR2X1 U14980 ( .A(n18230), .B(poly4_shifted[19]), .C(n17105), .D(n15823), 
        .Z(n15824) );
  COND1XL U14981 ( .A(n16775), .B(n18230), .C(n15824), .Z(n8854) );
  CANR2X1 U14982 ( .A(n12211), .B(Poly2[22]), .C(n16985), .D(poly2_shifted[22]), .Z(n15825) );
  COND1XL U14983 ( .A(n17001), .B(n12211), .C(n15825), .Z(n8988) );
  CANR2X1 U14984 ( .A(n12211), .B(Poly2[29]), .C(n16323), .D(poly2_shifted[29]), .Z(n15826) );
  COND1XL U14985 ( .A(n17185), .B(n12211), .C(n15826), .Z(n8981) );
  CIVX1 U14986 ( .A(n17742), .Z(n15827) );
  CANR2X1 U14987 ( .A(n12185), .B(poly11_shifted[15]), .C(n16323), .D(n15827), 
        .Z(n15828) );
  COND1XL U14988 ( .A(n17751), .B(n12185), .C(n15828), .Z(n11189) );
  CANR2X1 U14989 ( .A(n12211), .B(poly2_shifted[27]), .C(n17209), .D(
        poly2_shifted[15]), .Z(n15829) );
  COND1XL U14990 ( .A(n17196), .B(n12211), .C(n15829), .Z(n8995) );
  CANR2X1 U14991 ( .A(n12211), .B(Poly2[27]), .C(n16307), .D(poly2_shifted[27]), .Z(n15830) );
  COND1XL U14992 ( .A(n17741), .B(n12211), .C(n15830), .Z(n8983) );
  CANR2XL U14993 ( .A(n18198), .B(poly1_shifted[307]), .C(poly1_shifted[296]), 
        .D(n18017), .Z(n15831) );
  COND1XL U14994 ( .A(n17163), .B(n18198), .C(n15831), .Z(n9061) );
  CANR2X1 U14995 ( .A(n18198), .B(poly1_shifted[312]), .C(n17401), .D(
        poly1_shifted[301]), .Z(n15832) );
  COND1XL U14996 ( .A(n17090), .B(n18198), .C(n15832), .Z(n9056) );
  CANR2X1 U14997 ( .A(n17533), .B(poly0_shifted[189]), .C(n17314), .D(
        poly0_shifted[207]), .Z(n15833) );
  COND1XL U14998 ( .A(n17316), .B(n17185), .C(n15833), .Z(n9388) );
  CANR2X1 U14999 ( .A(n18234), .B(poly0_shifted[187]), .C(n17314), .D(
        poly0_shifted[205]), .Z(n15834) );
  COND1XL U15000 ( .A(n17316), .B(n17741), .C(n15834), .Z(n9390) );
  CANR2XL U15001 ( .A(n17574), .B(Poly7[235]), .C(n17285), .D(
        poly7_shifted[235]), .Z(n15835) );
  COND1XL U15002 ( .A(n16605), .B(n17574), .C(n15835), .Z(n9869) );
  CANR2X1 U15003 ( .A(n18230), .B(Poly4[30]), .C(n16502), .D(poly4_shifted[30]), .Z(n15836) );
  COND1XL U15004 ( .A(n17004), .B(n18230), .C(n15836), .Z(n8826) );
  CANR2X1 U15005 ( .A(n15737), .B(poly3_shifted[43]), .C(n17245), .D(
        poly3_shifted[29]), .Z(n15837) );
  COND1XL U15006 ( .A(n17185), .B(n15737), .C(n15837), .Z(n8911) );
  CENX1 U15007 ( .A(n17742), .B(Poly11[32]), .Z(n15838) );
  CANR2X1 U15008 ( .A(n17683), .B(Poly11[47]), .C(n17288), .D(n15838), .Z(
        n15839) );
  COND1XL U15009 ( .A(n17196), .B(n17747), .C(n15839), .Z(n11142) );
  CEOXL U15010 ( .A(Poly11[63]), .B(Poly11[84]), .Z(n15840) );
  CENX1 U15011 ( .A(n17742), .B(n15840), .Z(n15841) );
  CANR2X1 U15012 ( .A(n15843), .B(Poly11[78]), .C(n17198), .D(n15841), .Z(
        n15842) );
  COND1XL U15013 ( .A(n17699), .B(n15843), .C(n15842), .Z(n11111) );
  CENX1 U15014 ( .A(n15844), .B(Poly11[33]), .Z(n15845) );
  CANR2X1 U15015 ( .A(n17683), .B(Poly11[48]), .C(n17136), .D(n15845), .Z(
        n15846) );
  COND1XL U15016 ( .A(n17062), .B(n17747), .C(n15846), .Z(n11141) );
  CANR2X1 U15017 ( .A(n18230), .B(Poly4[22]), .C(n17334), .D(poly4_shifted[22]), .Z(n15847) );
  COND1XL U15018 ( .A(n17001), .B(n18230), .C(n15847), .Z(n8834) );
  CANR2X1 U15019 ( .A(n12211), .B(Poly2[24]), .C(n17458), .D(poly2_shifted[24]), .Z(n15848) );
  COND1XL U15020 ( .A(n17721), .B(n12211), .C(n15848), .Z(n8986) );
  CENX1 U15021 ( .A(n17680), .B(Poly11[34]), .Z(n15849) );
  CANR2X1 U15022 ( .A(n17683), .B(Poly11[49]), .C(n17527), .D(n15849), .Z(
        n15850) );
  COND1XL U15023 ( .A(n17076), .B(n17747), .C(n15850), .Z(n11140) );
  CANR2XL U15024 ( .A(n17411), .B(Poly10[41]), .C(n17206), .D(
        poly10_shifted[41]), .Z(n15851) );
  COND1XL U15025 ( .A(n17208), .B(n17411), .C(n15851), .Z(n11062) );
  CANR2X1 U15026 ( .A(n17731), .B(poly9_shifted[14]), .C(n17998), .D(
        Poly9[108]), .Z(n15852) );
  COND1XL U15027 ( .A(n13275), .B(n17731), .C(n15852), .Z(n11302) );
  CANR2X1 U15028 ( .A(n15737), .B(poly3_shifted[39]), .C(n17178), .D(
        poly3_shifted[25]), .Z(n15853) );
  COND1XL U15029 ( .A(n17123), .B(n15737), .C(n15853), .Z(n8915) );
  CIVXL U15030 ( .A(n17692), .Z(n15854) );
  CANR2X1 U15031 ( .A(n12211), .B(poly2_shifted[14]), .C(n17375), .D(n15854), 
        .Z(n15855) );
  COND1XL U15032 ( .A(n16775), .B(n12211), .C(n15855), .Z(n9008) );
  CEOXL U15033 ( .A(Poly8[95]), .B(Poly8[16]), .Z(n15856) );
  CANR2X1 U15034 ( .A(n12175), .B(poly8_shifted[44]), .C(n17203), .D(n15856), 
        .Z(n15857) );
  COND1XL U15035 ( .A(n13418), .B(n12175), .C(n15857), .Z(n11371) );
  CANR2X1 U15036 ( .A(n12211), .B(poly2_shifted[18]), .C(n17105), .D(Poly2[64]), .Z(n15858) );
  COND1XL U15037 ( .A(n17757), .B(n12211), .C(n15858), .Z(n9004) );
  CENX1 U15038 ( .A(Poly11[46]), .B(n15859), .Z(n15860) );
  CANR2X1 U15039 ( .A(n17747), .B(Poly11[61]), .C(n17099), .D(n15860), .Z(
        n15861) );
  COND1XL U15040 ( .A(n17185), .B(n17747), .C(n15861), .Z(n11128) );
  CIVXL U15041 ( .A(n15971), .Z(n15862) );
  CANR2X1 U15042 ( .A(n12211), .B(poly2_shifted[12]), .C(n16307), .D(n15862), 
        .Z(n15863) );
  COND1XL U15043 ( .A(n17751), .B(n12211), .C(n15863), .Z(n9010) );
  CANR2X1 U15044 ( .A(n18230), .B(Poly4[16]), .C(n16502), .D(Poly4[60]), .Z(
        n15864) );
  COND1XL U15045 ( .A(n17062), .B(n18230), .C(n15864), .Z(n8840) );
  CANR2X1 U15046 ( .A(poly4_shifted[17]), .B(n18230), .C(n16787), .D(n15865), 
        .Z(n15866) );
  COND1XL U15047 ( .A(n17751), .B(n18230), .C(n15866), .Z(n8856) );
  CANR2X1 U15048 ( .A(n17053), .B(Poly1[202]), .C(n16312), .D(
        poly1_shifted[202]), .Z(n15867) );
  COND1XL U15049 ( .A(n12014), .B(n17053), .C(n15867), .Z(n9155) );
  CANR2X1 U15050 ( .A(n12153), .B(Poly4[32]), .C(n16502), .D(poly4_shifted[32]), .Z(n15868) );
  COND1XL U15051 ( .A(n17751), .B(n12153), .C(n15868), .Z(n8824) );
  CANR2X1 U15052 ( .A(n17750), .B(Poly8[67]), .C(n16323), .D(poly8_shifted[67]), .Z(n15869) );
  COND1XL U15053 ( .A(n13275), .B(n17750), .C(n15869), .Z(n11334) );
  CANR2X1 U15054 ( .A(n12192), .B(Poly1[226]), .C(n16488), .D(
        poly1_shifted[226]), .Z(n15870) );
  COND1XL U15055 ( .A(n16775), .B(n12192), .C(n15870), .Z(n9131) );
  CENX1 U15056 ( .A(Poly8[89]), .B(Poly8[91]), .Z(n15871) );
  CENX1 U15057 ( .A(Poly8[10]), .B(n15871), .Z(n15872) );
  CANR2X1 U15058 ( .A(n12175), .B(poly8_shifted[38]), .C(n16323), .D(n15872), 
        .Z(n15873) );
  COND1XL U15059 ( .A(n17721), .B(n12175), .C(n15873), .Z(n11377) );
  CEOXL U15060 ( .A(Poly10[42]), .B(Poly10[26]), .Z(n15874) );
  CANR2X1 U15061 ( .A(n17411), .B(Poly10[38]), .C(n17523), .D(n15874), .Z(
        n15875) );
  COND1XL U15062 ( .A(n16779), .B(n17411), .C(n15875), .Z(n11065) );
  CANR2X1 U15063 ( .A(n12211), .B(poly2_shifted[20]), .C(n16323), .D(Poly2[66]), .Z(n15876) );
  COND1XL U15064 ( .A(n17163), .B(n12211), .C(n15876), .Z(n9002) );
  CANR2X1 U15065 ( .A(n18230), .B(Poly4[17]), .C(n16502), .D(poly4_shifted[17]), .Z(n15877) );
  COND1XL U15066 ( .A(n17173), .B(n18230), .C(n15877), .Z(n8839) );
  CANR2X1 U15067 ( .A(n18230), .B(Poly4[24]), .C(n17334), .D(poly4_shifted[24]), .Z(n15878) );
  COND1XL U15068 ( .A(n17721), .B(n18230), .C(n15878), .Z(n8832) );
  CENX1 U15069 ( .A(Poly0[104]), .B(Poly0[203]), .Z(n15879) );
  COND1XL U15070 ( .A(n15879), .B(n17959), .C(n13367), .Z(n15881) );
  CMX2XL U15071 ( .A0(n15881), .A1(poly0_shifted[140]), .S(n15880), .Z(n9455)
         );
  CANR2X1 U15072 ( .A(n13351), .B(poly9_shifted[59]), .C(n16702), .D(
        poly9_shifted[48]), .Z(n15882) );
  COND1XL U15073 ( .A(n17062), .B(n13351), .C(n15882), .Z(n11257) );
  CANR2X1 U15074 ( .A(n13351), .B(poly9_shifted[52]), .C(n16919), .D(
        poly9_shifted[41]), .Z(n15883) );
  COND1XL U15075 ( .A(n12002), .B(n13351), .C(n15883), .Z(n11264) );
  CANR2X1 U15076 ( .A(n13351), .B(poly9_shifted[67]), .C(n16372), .D(
        poly9_shifted[56]), .Z(n15884) );
  COND1XL U15077 ( .A(n17721), .B(n13351), .C(n15884), .Z(n11249) );
  CANR2X1 U15078 ( .A(n13351), .B(poly9_shifted[54]), .C(n18234), .D(
        poly9_shifted[43]), .Z(n15885) );
  COND1XL U15079 ( .A(n16605), .B(n13351), .C(n15885), .Z(n11262) );
  CANR2X1 U15080 ( .A(n13351), .B(poly9_shifted[53]), .C(n17362), .D(
        poly9_shifted[42]), .Z(n15886) );
  COND1XL U15081 ( .A(n12014), .B(n13351), .C(n15886), .Z(n11263) );
  CANR2X1 U15082 ( .A(n13351), .B(poly9_shifted[68]), .C(n17705), .D(
        poly9_shifted[57]), .Z(n15887) );
  COND1XL U15083 ( .A(n17200), .B(n13351), .C(n15887), .Z(n11248) );
  CANR2X1 U15084 ( .A(n13351), .B(poly9_shifted[72]), .C(n17705), .D(
        poly9_shifted[61]), .Z(n15888) );
  COND1XL U15085 ( .A(n17185), .B(n13351), .C(n15888), .Z(n11244) );
  CEOXL U15086 ( .A(Poly9[115]), .B(Poly9[26]), .Z(n15889) );
  CANR2X1 U15087 ( .A(n13351), .B(poly9_shifted[48]), .C(n16644), .D(n15889), 
        .Z(n15890) );
  COND1XL U15088 ( .A(n11981), .B(n13351), .C(n15890), .Z(n11268) );
  CANR2XL U15089 ( .A(n13351), .B(poly9_shifted[70]), .C(poly9_shifted[59]), 
        .D(n18017), .Z(n15891) );
  COND1XL U15090 ( .A(n17741), .B(n13351), .C(n15891), .Z(n11246) );
  CANR2X1 U15091 ( .A(n13351), .B(poly9_shifted[51]), .C(n17466), .D(
        poly9_shifted[40]), .Z(n15892) );
  COND1XL U15092 ( .A(n17163), .B(n13351), .C(n15892), .Z(n11265) );
  CANR2X1 U15093 ( .A(n13351), .B(poly9_shifted[56]), .C(n17714), .D(
        poly9_shifted[45]), .Z(n15893) );
  COND1XL U15094 ( .A(n17090), .B(n13351), .C(n15893), .Z(n11260) );
  CANR2X1 U15095 ( .A(n18230), .B(Poly4[27]), .C(n17295), .D(poly4_shifted[27]), .Z(n15894) );
  COND1XL U15096 ( .A(n17741), .B(n18230), .C(n15894), .Z(n8829) );
  CANR2X1 U15097 ( .A(n18198), .B(poly1_shifted[306]), .C(n17655), .D(
        poly1_shifted[295]), .Z(n15895) );
  COND1XL U15098 ( .A(n17718), .B(n18198), .C(n15895), .Z(n9062) );
  CANR2X1 U15099 ( .A(n18198), .B(poly1_shifted[309]), .C(n17642), .D(
        poly1_shifted[298]), .Z(n15896) );
  COND1XL U15100 ( .A(n12014), .B(n18198), .C(n15896), .Z(n9059) );
  CANR2X1 U15101 ( .A(n18198), .B(poly1_shifted[304]), .C(n17705), .D(
        poly1_shifted[293]), .Z(n15897) );
  COND1XL U15102 ( .A(n11983), .B(n18198), .C(n15897), .Z(n9064) );
  CANR2XL U15103 ( .A(n17430), .B(Poly13[519]), .C(n17607), .D(
        poly13_shifted[519]), .Z(n15898) );
  COND1XL U15104 ( .A(n16939), .B(n17430), .C(n15898), .Z(n10541) );
  CANR2X1 U15105 ( .A(n12900), .B(poly13_shifted[49]), .C(n17072), .D(
        poly13_shifted[35]), .Z(n15899) );
  COND1XL U15106 ( .A(n13275), .B(n12900), .C(n15899), .Z(n11025) );
  CANR2X1 U15107 ( .A(n12900), .B(poly13_shifted[76]), .C(n17266), .D(
        poly13_shifted[62]), .Z(n15900) );
  COND1XL U15108 ( .A(n13418), .B(n12900), .C(n15900), .Z(n10998) );
  CANR2X1 U15109 ( .A(n12900), .B(poly13_shifted[61]), .C(n17401), .D(
        poly13_shifted[47]), .Z(n15901) );
  COND1XL U15110 ( .A(n17196), .B(n12900), .C(n15901), .Z(n11013) );
  CANR2X1 U15111 ( .A(n12900), .B(poly13_shifted[62]), .C(n17266), .D(
        poly13_shifted[48]), .Z(n15902) );
  COND1XL U15112 ( .A(n17062), .B(n12900), .C(n15902), .Z(n11012) );
  CANR2X1 U15113 ( .A(n12900), .B(poly13_shifted[48]), .C(n17266), .D(
        poly13_shifted[34]), .Z(n15903) );
  COND1XL U15114 ( .A(n16775), .B(n12900), .C(n15903), .Z(n11026) );
  CMXI2XL U15115 ( .A0(n18138), .A1(poly10_shifted[19]), .S(n17962), .Z(n15904) );
  COND1XL U15116 ( .A(n17495), .B(n15905), .C(n15904), .Z(n11096) );
  CANR2X1 U15117 ( .A(n12008), .B(poly14_shifted[166]), .C(n17714), .D(
        poly14_shifted[150]), .Z(n15906) );
  COND1XL U15118 ( .A(n17001), .B(n12008), .C(n15906), .Z(n10255) );
  CIVX1 U15119 ( .A(Poly5[78]), .Z(n17939) );
  CANR2X1 U15120 ( .A(n17045), .B(n18160), .C(n17158), .D(poly5_shifted[78]), 
        .Z(n15907) );
  COND1XL U15121 ( .A(n17045), .B(n17939), .C(n15907), .Z(n11448) );
  CANR2X1 U15122 ( .A(n17955), .B(poly9_shifted[88]), .C(n16427), .D(
        poly9_shifted[77]), .Z(n15908) );
  COND1XL U15123 ( .A(n17065), .B(n17955), .C(n15908), .Z(n11228) );
  CANR2X1 U15124 ( .A(n17955), .B(poly9_shifted[87]), .C(n18047), .D(
        poly9_shifted[76]), .Z(n15909) );
  COND1XL U15125 ( .A(n17218), .B(n17955), .C(n15909), .Z(n11229) );
  CANR2X1 U15126 ( .A(n17955), .B(Poly9[94]), .C(n17458), .D(poly9_shifted[94]), .Z(n15910) );
  COND1XL U15127 ( .A(n13418), .B(n17955), .C(n15910), .Z(n11211) );
  CANR2X1 U15128 ( .A(n17955), .B(Poly9[92]), .C(n17538), .D(poly9_shifted[92]), .Z(n15911) );
  COND1XL U15129 ( .A(n11978), .B(n17955), .C(n15911), .Z(n11213) );
  CANR2XL U15130 ( .A(n17955), .B(Poly9[86]), .C(poly9_shifted[86]), .D(n18017), .Z(n15912) );
  COND1XL U15131 ( .A(n17753), .B(n17955), .C(n15912), .Z(n11219) );
  CANR2X1 U15132 ( .A(n17955), .B(poly9_shifted[91]), .C(n17105), .D(
        poly9_shifted[80]), .Z(n15913) );
  COND1XL U15133 ( .A(n17062), .B(n17955), .C(n15913), .Z(n11225) );
  CANR2X1 U15134 ( .A(n17491), .B(poly13_shifted[494]), .C(n17634), .D(
        poly13_shifted[480]), .Z(n15914) );
  COND1XL U15135 ( .A(n17751), .B(n17491), .C(n15914), .Z(n10580) );
  CANR2X1 U15136 ( .A(n17491), .B(poly13_shifted[510]), .C(n17755), .D(
        poly13_shifted[496]), .Z(n15915) );
  COND1XL U15137 ( .A(n17062), .B(n17491), .C(n15915), .Z(n10564) );
  CAN2XL U15138 ( .A(n18017), .B(Poly12[126]), .Z(n15916) );
  CANR1XL U15139 ( .A(Poly12[15]), .B(n12997), .C(n15916), .Z(n15917) );
  COND1XL U15140 ( .A(n17196), .B(n12997), .C(n15917), .Z(n10517) );
  CEOXL U15141 ( .A(Poly7[405]), .B(dataselector[62]), .Z(n15918) );
  CENX1 U15142 ( .A(n15919), .B(n15918), .Z(n15921) );
  CANR2X1 U15143 ( .A(n14716), .B(n17832), .C(dataselector[1]), .D(n16410), 
        .Z(n15920) );
  COND1XL U15144 ( .A(n17829), .B(n15921), .C(n15920), .Z(n8794) );
  CANR2X1 U15145 ( .A(n17376), .B(Poly15[56]), .C(n16540), .D(
        poly15_shifted[56]), .Z(n15922) );
  COND1XL U15146 ( .A(n17721), .B(n17376), .C(n15922), .Z(n9581) );
  CANR2X1 U15147 ( .A(n18230), .B(Poly4[31]), .C(n17334), .D(poly4_shifted[31]), .Z(n15923) );
  COND1XL U15148 ( .A(n17188), .B(n18230), .C(n15923), .Z(n8825) );
  CANR2X1 U15149 ( .A(n12210), .B(poly1_shifted[202]), .C(n16312), .D(
        poly1_shifted[191]), .Z(n15924) );
  COND1XL U15150 ( .A(n17188), .B(n12210), .C(n15924), .Z(n9166) );
  CEOXL U15151 ( .A(Poly2[51]), .B(n15971), .Z(n15925) );
  CENX1 U15152 ( .A(Poly2[63]), .B(n15925), .Z(n15926) );
  CANR2X1 U15153 ( .A(n17306), .B(Poly2[63]), .C(n16479), .D(n15926), .Z(
        n15927) );
  COND1XL U15154 ( .A(n17188), .B(n17306), .C(n15927), .Z(n8947) );
  CANR2X1 U15155 ( .A(n17053), .B(poly1_shifted[234]), .C(n16479), .D(
        poly1_shifted[223]), .Z(n15928) );
  COND1XL U15156 ( .A(n17188), .B(n17053), .C(n15928), .Z(n9134) );
  CANR2X1 U15157 ( .A(n12598), .B(Poly12[63]), .C(n18234), .D(
        poly12_shifted[63]), .Z(n15929) );
  COND1XL U15158 ( .A(n17188), .B(n12598), .C(n15929), .Z(n10469) );
  CANR2XL U15159 ( .A(n18198), .B(poly1_shifted[330]), .C(poly1_shifted[319]), 
        .D(n18017), .Z(n15930) );
  COND1XL U15160 ( .A(n17188), .B(n18198), .C(n15930), .Z(n9038) );
  CANR2X1 U15161 ( .A(n12932), .B(Poly14[287]), .C(n17523), .D(
        poly14_shifted[287]), .Z(n15931) );
  COND1XL U15162 ( .A(n17188), .B(n12932), .C(n15931), .Z(n10118) );
  CANR2X1 U15163 ( .A(n12012), .B(poly1_shifted[106]), .C(n17203), .D(
        poly1_shifted[95]), .Z(n15932) );
  COND1XL U15164 ( .A(n17188), .B(n12012), .C(n15932), .Z(n9262) );
  CANR2X1 U15165 ( .A(n12009), .B(poly14_shifted[143]), .C(n17535), .D(
        poly14_shifted[127]), .Z(n15933) );
  COND1XL U15166 ( .A(n17188), .B(n12009), .C(n15933), .Z(n10278) );
  CANR2X1 U15167 ( .A(n15737), .B(Poly3[31]), .C(n17158), .D(poly3_shifted[31]), .Z(n15934) );
  COND1XL U15168 ( .A(n17188), .B(n15737), .C(n15934), .Z(n8909) );
  CANR2X1 U15169 ( .A(n12008), .B(poly14_shifted[175]), .C(n17362), .D(
        poly14_shifted[159]), .Z(n15935) );
  COND1XL U15170 ( .A(n17188), .B(n12008), .C(n15935), .Z(n10246) );
  CANR2X1 U15171 ( .A(n17444), .B(Poly14[297]), .C(n17266), .D(
        poly14_shifted[297]), .Z(n15936) );
  COND1XL U15172 ( .A(n17208), .B(n17444), .C(n15936), .Z(n10108) );
  CANR2X1 U15173 ( .A(n17444), .B(Poly14[293]), .C(n16435), .D(
        poly14_shifted[293]), .Z(n15937) );
  COND1XL U15174 ( .A(n11991), .B(n17444), .C(n15937), .Z(n10112) );
  CANR2X1 U15175 ( .A(n17444), .B(Poly14[299]), .C(n16307), .D(
        poly14_shifted[299]), .Z(n15938) );
  COND1XL U15176 ( .A(n16605), .B(n17444), .C(n15938), .Z(n10106) );
  CANR2X1 U15177 ( .A(n17444), .B(Poly14[291]), .C(n17714), .D(
        poly14_shifted[291]), .Z(n15939) );
  COND1XL U15178 ( .A(n13275), .B(n17444), .C(n15939), .Z(n10114) );
  CMXI2XL U15179 ( .A0(n18142), .A1(poly10_shifted[20]), .S(n17962), .Z(n15940) );
  COND1XL U15180 ( .A(n15941), .B(n17495), .C(n15940), .Z(n11095) );
  CIVX1 U15181 ( .A(n15942), .Z(n15944) );
  CMXI2X1 U15182 ( .A0(n14754), .A1(poly10_shifted[18]), .S(n17962), .Z(n15943) );
  COND1XL U15183 ( .A(n17959), .B(n15944), .C(n15943), .Z(n11097) );
  CMXI2XL U15184 ( .A0(n16381), .A1(Poly10[11]), .S(n17962), .Z(n15945) );
  COND1XL U15185 ( .A(n15946), .B(n17959), .C(n15945), .Z(n11092) );
  CMXI2XL U15186 ( .A0(n18189), .A1(poly10_shifted[21]), .S(n17962), .Z(n15947) );
  COND1XL U15187 ( .A(n15948), .B(n17829), .C(n15947), .Z(n11094) );
  CIVXL U15188 ( .A(Poly10[31]), .Z(n15950) );
  CMXI2XL U15189 ( .A0(n18108), .A1(Poly10[0]), .S(n17962), .Z(n15949) );
  COND1XL U15190 ( .A(n15950), .B(n17959), .C(n15949), .Z(n11103) );
  CIVXL U15191 ( .A(n15951), .Z(n15953) );
  CMXI2X1 U15192 ( .A0(n11990), .A1(poly10_shifted[17]), .S(n17962), .Z(n15952) );
  COND1XL U15193 ( .A(n17959), .B(n15953), .C(n15952), .Z(n11098) );
  CMXI2X1 U15194 ( .A0(n18053), .A1(Poly10[3]), .S(n17962), .Z(n15954) );
  COND1XL U15195 ( .A(n17744), .B(n15955), .C(n15954), .Z(n11100) );
  CANR2X1 U15196 ( .A(n12161), .B(Poly12[94]), .C(n16985), .D(
        poly12_shifted[94]), .Z(n15956) );
  COND1XL U15197 ( .A(n13418), .B(n12161), .C(n15956), .Z(n10438) );
  CANR2X1 U15198 ( .A(n12161), .B(Poly12[91]), .C(n16488), .D(
        poly12_shifted[91]), .Z(n15957) );
  COND1XL U15199 ( .A(n17741), .B(n12161), .C(n15957), .Z(n10441) );
  CANR2X1 U15200 ( .A(n12161), .B(Poly12[86]), .C(n17705), .D(
        poly12_shifted[86]), .Z(n15958) );
  COND1XL U15201 ( .A(n17001), .B(n12161), .C(n15958), .Z(n10446) );
  CANR2X1 U15202 ( .A(n12900), .B(poly13_shifted[74]), .C(n18234), .D(
        poly13_shifted[60]), .Z(n15959) );
  COND1XL U15203 ( .A(n11978), .B(n12900), .C(n15959), .Z(n11000) );
  CENX1 U15204 ( .A(Poly0[157]), .B(Poly0[209]), .Z(n15962) );
  COND2X1 U15205 ( .A(n15960), .B(poly0_shifted[193]), .C(n18206), .D(n17314), 
        .Z(n15961) );
  COND1XL U15206 ( .A(n15962), .B(n17744), .C(n15961), .Z(n9402) );
  CANR2X1 U15207 ( .A(n17430), .B(Poly13[523]), .C(n17668), .D(
        poly13_shifted[523]), .Z(n15963) );
  COND1XL U15208 ( .A(n16994), .B(n17430), .C(n15963), .Z(n10537) );
  CANR2X1 U15209 ( .A(n12262), .B(Poly9[107]), .C(n17209), .D(
        poly9_shifted[107]), .Z(n15964) );
  COND1XL U15210 ( .A(n16994), .B(n12262), .C(n15964), .Z(n11198) );
  CANR2X1 U15211 ( .A(n12958), .B(poly14_shifted[91]), .C(n17063), .D(
        poly14_shifted[75]), .Z(n15965) );
  COND1XL U15212 ( .A(n16994), .B(n12958), .C(n15965), .Z(n10330) );
  CAN2XL U15213 ( .A(n18017), .B(Poly13[525]), .Z(n15966) );
  CANR1XL U15214 ( .A(poly13_shifted[25]), .B(n13124), .C(n15966), .Z(n15967)
         );
  COND1XL U15215 ( .A(n16994), .B(n13124), .C(n15967), .Z(n11049) );
  CANR2X1 U15216 ( .A(n12009), .B(poly14_shifted[123]), .C(n17063), .D(
        poly14_shifted[107]), .Z(n15968) );
  COND1XL U15217 ( .A(n16994), .B(n12009), .C(n15968), .Z(n10298) );
  CANR2X1 U15218 ( .A(n12012), .B(poly1_shifted[86]), .C(n16479), .D(
        poly1_shifted[75]), .Z(n15969) );
  COND1XL U15219 ( .A(n16994), .B(n12012), .C(n15969), .Z(n9282) );
  CENX1 U15220 ( .A(Poly2[31]), .B(Poly2[67]), .Z(n15970) );
  CENX1 U15221 ( .A(n15971), .B(n15970), .Z(n15972) );
  CNR2X1 U15222 ( .A(n15972), .B(n15673), .Z(n15973) );
  CANR1XL U15223 ( .A(poly2_shifted[55]), .B(n17306), .C(n15973), .Z(n15974)
         );
  COND1XL U15224 ( .A(n16994), .B(n17306), .C(n15974), .Z(n8967) );
  CANR2X1 U15225 ( .A(n17043), .B(Poly13[395]), .C(n17072), .D(
        poly13_shifted[395]), .Z(n15975) );
  COND1XL U15226 ( .A(n16994), .B(n17043), .C(n15975), .Z(n10665) );
  CEOXL U15227 ( .A(Poly7[401]), .B(Poly7[406]), .Z(n15976) );
  CENX1 U15228 ( .A(Poly7[185]), .B(n15976), .Z(n15977) );
  CNR2XL U15229 ( .A(n15977), .B(n17829), .Z(n15978) );
  CANR1XL U15230 ( .A(poly7_shifted[209]), .B(n17273), .C(n15978), .Z(n15979)
         );
  COND1XL U15231 ( .A(n11993), .B(n17273), .C(n15979), .Z(n9907) );
  CENX1 U15232 ( .A(dataselector[59]), .B(dataselector[51]), .Z(n15980) );
  CENX1 U15233 ( .A(n15981), .B(n15980), .Z(n15983) );
  CANR2X1 U15234 ( .A(n18095), .B(n18248), .C(n16350), .D(dataselector[58]), 
        .Z(n15982) );
  COND1XL U15235 ( .A(n17959), .B(n15983), .C(n15982), .Z(n8737) );
  CANR2X1 U15236 ( .A(n13124), .B(poly13_shifted[14]), .C(n17705), .D(
        Poly13[514]), .Z(n15984) );
  COND1XL U15237 ( .A(n12011), .B(n13124), .C(n15984), .Z(n11060) );
  CANR2XL U15238 ( .A(n12932), .B(poly14_shifted[272]), .C(poly14_shifted[256]), .D(n18017), .Z(n15985) );
  COND1XL U15239 ( .A(n12011), .B(n12932), .C(n15985), .Z(n10149) );
  CANR2XL U15240 ( .A(n17667), .B(poly13_shifted[206]), .C(n17755), .D(
        poly13_shifted[192]), .Z(n15986) );
  COND1XL U15241 ( .A(n12011), .B(n17667), .C(n15986), .Z(n10868) );
  CANR2XL U15242 ( .A(n17444), .B(Poly14[288]), .C(n18234), .D(
        poly14_shifted[288]), .Z(n15987) );
  COND1XL U15243 ( .A(n12011), .B(n17444), .C(n15987), .Z(n10117) );
  CANR2X1 U15244 ( .A(n13129), .B(poly14_shifted[176]), .C(n17755), .D(
        poly14_shifted[160]), .Z(n15988) );
  COND1XL U15245 ( .A(n12011), .B(n13129), .C(n15988), .Z(n10245) );
  CANR2X1 U15246 ( .A(n12008), .B(poly14_shifted[144]), .C(n17535), .D(
        poly14_shifted[128]), .Z(n15989) );
  COND1XL U15247 ( .A(n12011), .B(n12008), .C(n15989), .Z(n10277) );
  CANR2X1 U15248 ( .A(n17731), .B(poly9_shifted[11]), .C(n17755), .D(
        Poly9[105]), .Z(n15990) );
  COND1XL U15249 ( .A(n12011), .B(n17731), .C(n15990), .Z(n11305) );
  CANR2X1 U15250 ( .A(n17430), .B(poly13_shifted[526]), .C(n17362), .D(
        poly13_shifted[512]), .Z(n15991) );
  COND1XL U15251 ( .A(n12011), .B(n17430), .C(n15991), .Z(n10548) );
  CAN2XL U15252 ( .A(n18017), .B(poly13_shifted[32]), .Z(n15992) );
  CANR1XL U15253 ( .A(poly13_shifted[46]), .B(n12900), .C(n15992), .Z(n15993)
         );
  COND1XL U15254 ( .A(n12011), .B(n12900), .C(n15993), .Z(n11028) );
  CANR2XL U15255 ( .A(n17942), .B(poly5_shifted[78]), .C(n16326), .D(
        poly5_shifted[64]), .Z(n15994) );
  COND1XL U15256 ( .A(n12011), .B(n17942), .C(n15994), .Z(n11462) );
  CANR2X1 U15257 ( .A(n12009), .B(poly14_shifted[112]), .C(n17401), .D(
        poly14_shifted[96]), .Z(n15995) );
  COND1XL U15258 ( .A(n12011), .B(n12009), .C(n15995), .Z(n10309) );
  CEOXL U15259 ( .A(Poly4[32]), .B(Poly4[46]), .Z(n15996) );
  CENX1 U15260 ( .A(n16988), .B(n15996), .Z(n15998) );
  CMXI2XL U15261 ( .A0(n14297), .A1(Poly4[49]), .S(n12153), .Z(n15997) );
  COND1XL U15262 ( .A(n15998), .B(n17829), .C(n15997), .Z(n8807) );
  CANR2X1 U15263 ( .A(n12977), .B(Poly7[184]), .C(n17535), .D(
        poly7_shifted[184]), .Z(n15999) );
  COND1XL U15264 ( .A(n17721), .B(n12977), .C(n15999), .Z(n9920) );
  CANR2X1 U15265 ( .A(n12977), .B(Poly7[185]), .C(n17533), .D(
        poly7_shifted[185]), .Z(n16000) );
  COND1XL U15266 ( .A(n17200), .B(n12977), .C(n16000), .Z(n9919) );
  CANR2X1 U15267 ( .A(n12977), .B(poly7_shifted[172]), .C(n17209), .D(
        poly7_shifted[160]), .Z(n16001) );
  COND1XL U15268 ( .A(n12011), .B(n12977), .C(n16001), .Z(n9944) );
  CANR2X1 U15269 ( .A(n12977), .B(poly7_shifted[181]), .C(n17178), .D(
        poly7_shifted[169]), .Z(n16002) );
  COND1XL U15270 ( .A(n17208), .B(n12977), .C(n16002), .Z(n9935) );
  CANR2X1 U15271 ( .A(n12977), .B(poly7_shifted[177]), .C(n16479), .D(
        poly7_shifted[165]), .Z(n16003) );
  COND1XL U15272 ( .A(n11983), .B(n12977), .C(n16003), .Z(n9939) );
  CANR2X1 U15273 ( .A(n12977), .B(poly7_shifted[185]), .C(n17533), .D(
        poly7_shifted[173]), .Z(n16004) );
  COND1XL U15274 ( .A(n17090), .B(n12977), .C(n16004), .Z(n9931) );
  CANR2X1 U15275 ( .A(n17045), .B(n18082), .C(n17755), .D(poly5_shifted[84]), 
        .Z(n16005) );
  COND1XL U15276 ( .A(n17045), .B(n16006), .C(n16005), .Z(n11442) );
  CAN2XL U15277 ( .A(n18017), .B(poly14_shifted[39]), .Z(n16007) );
  CANR1XL U15278 ( .A(poly14_shifted[55]), .B(n17525), .C(n16007), .Z(n16008)
         );
  COND1XL U15279 ( .A(n16939), .B(n17525), .C(n16008), .Z(n10366) );
  CANR2X1 U15280 ( .A(n13124), .B(poly13_shifted[43]), .C(n17508), .D(
        poly13_shifted[29]), .Z(n16009) );
  COND1XL U15281 ( .A(n17185), .B(n13124), .C(n16009), .Z(n11031) );
  CANR2X1 U15282 ( .A(n13124), .B(poly13_shifted[17]), .C(n17620), .D(
        Poly13[517]), .Z(n16010) );
  COND1XL U15283 ( .A(n13275), .B(n13124), .C(n16010), .Z(n11057) );
  CANR2X1 U15284 ( .A(n13124), .B(poly13_shifted[23]), .C(n17668), .D(
        Poly13[523]), .Z(n16011) );
  COND1XL U15285 ( .A(n17208), .B(n13124), .C(n16011), .Z(n11051) );
  CANR2X1 U15286 ( .A(n17750), .B(Poly8[95]), .C(n17398), .D(poly8_shifted[95]), .Z(n16012) );
  COND1XL U15287 ( .A(n17188), .B(n17750), .C(n16012), .Z(n11306) );
  CANR2X1 U15288 ( .A(n12161), .B(Poly12[95]), .C(n18234), .D(
        poly12_shifted[95]), .Z(n16013) );
  COND1XL U15289 ( .A(n17188), .B(n12161), .C(n16013), .Z(n10437) );
  CANR2X1 U15290 ( .A(n12900), .B(poly13_shifted[66]), .C(n17094), .D(
        poly13_shifted[52]), .Z(n16014) );
  COND1XL U15291 ( .A(n17707), .B(n12900), .C(n16014), .Z(n11008) );
  CANR2X1 U15292 ( .A(n13124), .B(poly13_shifted[24]), .C(n17295), .D(
        Poly13[524]), .Z(n16015) );
  COND1XL U15293 ( .A(n12014), .B(n13124), .C(n16015), .Z(n11050) );
  CANR2X1 U15294 ( .A(n12900), .B(poly13_shifted[58]), .C(n17466), .D(
        poly13_shifted[44]), .Z(n16016) );
  COND1XL U15295 ( .A(n17087), .B(n12900), .C(n16016), .Z(n11016) );
  CEOXL U15296 ( .A(Poly13[524]), .B(Poly13[279]), .Z(n16017) );
  CANR2X1 U15297 ( .A(n17615), .B(poly13_shifted[307]), .C(n17613), .D(n16017), 
        .Z(n16018) );
  COND1XL U15298 ( .A(n11993), .B(n17615), .C(n16018), .Z(n10767) );
  CANR2X1 U15299 ( .A(n13124), .B(poly13_shifted[38]), .C(n16583), .D(
        poly13_shifted[24]), .Z(n16019) );
  COND1XL U15300 ( .A(n17721), .B(n13124), .C(n16019), .Z(n11036) );
  CANR2X1 U15301 ( .A(n16425), .B(poly1_shifted[136]), .C(n17466), .D(
        poly1_shifted[125]), .Z(n16020) );
  COND1XL U15302 ( .A(n17185), .B(n16425), .C(n16020), .Z(n9232) );
  CANR2X1 U15303 ( .A(n16425), .B(poly1_shifted[129]), .C(n17266), .D(
        poly1_shifted[118]), .Z(n16021) );
  COND1XL U15304 ( .A(n17001), .B(n16425), .C(n16021), .Z(n9239) );
  CANR2X1 U15305 ( .A(n18002), .B(poly14_shifted[25]), .C(n17362), .D(
        Poly14[294]), .Z(n16022) );
  COND1XL U15306 ( .A(n17208), .B(n18002), .C(n16022), .Z(n10396) );
  CANR2X1 U15307 ( .A(n12009), .B(poly14_shifted[121]), .C(n17362), .D(
        poly14_shifted[105]), .Z(n16023) );
  COND1XL U15308 ( .A(n17208), .B(n12009), .C(n16023), .Z(n10300) );
  CANR2X1 U15309 ( .A(n17444), .B(Poly14[290]), .C(n16427), .D(
        poly14_shifted[290]), .Z(n16024) );
  COND1XL U15310 ( .A(n16303), .B(n17444), .C(n16024), .Z(n10115) );
  CANR2X1 U15311 ( .A(n12932), .B(poly14_shifted[274]), .C(n17504), .D(
        poly14_shifted[258]), .Z(n16025) );
  COND1XL U15312 ( .A(n16303), .B(n12932), .C(n16025), .Z(n10147) );
  CANR2X1 U15313 ( .A(n18002), .B(poly14_shifted[31]), .C(n17965), .D(
        Poly14[300]), .Z(n16026) );
  COND1XL U15314 ( .A(n17196), .B(n18002), .C(n16026), .Z(n10390) );
  CANR2X1 U15315 ( .A(n17444), .B(Poly14[298]), .C(n17362), .D(
        poly14_shifted[298]), .Z(n16027) );
  COND1XL U15316 ( .A(n12014), .B(n17444), .C(n16027), .Z(n10107) );
  CANR2X1 U15317 ( .A(n17935), .B(poly5_shifted[74]), .C(n17266), .D(
        poly5_shifted[60]), .Z(n16028) );
  COND1XL U15318 ( .A(n11978), .B(n17935), .C(n16028), .Z(n11466) );
  CANR2X1 U15319 ( .A(n18002), .B(poly14_shifted[37]), .C(n17998), .D(
        poly14_shifted[21]), .Z(n16029) );
  COND1XL U15320 ( .A(n12006), .B(n18002), .C(n16029), .Z(n10384) );
  CANR2X1 U15321 ( .A(n16425), .B(poly1_shifted[116]), .C(n17533), .D(
        poly1_shifted[105]), .Z(n16030) );
  COND1XL U15322 ( .A(n17208), .B(n16425), .C(n16030), .Z(n9252) );
  CANR2X1 U15323 ( .A(n17053), .B(Poly1[203]), .C(n17121), .D(
        poly1_shifted[203]), .Z(n16031) );
  COND1XL U15324 ( .A(n16605), .B(n17053), .C(n16031), .Z(n9154) );
  CANR2X1 U15325 ( .A(n12008), .B(poly14_shifted[155]), .C(n17063), .D(
        poly14_shifted[139]), .Z(n16032) );
  COND1XL U15326 ( .A(n16605), .B(n12008), .C(n16032), .Z(n10266) );
  CANR2X1 U15327 ( .A(n17750), .B(Poly8[75]), .C(n16307), .D(poly8_shifted[75]), .Z(n16033) );
  COND1XL U15328 ( .A(n16605), .B(n17750), .C(n16033), .Z(n11326) );
  CANR2X1 U15329 ( .A(n12997), .B(Poly12[29]), .C(n17640), .D(
        poly12_shifted[29]), .Z(n16034) );
  COND1XL U15330 ( .A(n17185), .B(n12997), .C(n16034), .Z(n10503) );
  CANR2X1 U15331 ( .A(n12997), .B(Poly12[17]), .C(n17238), .D(
        poly12_shifted[17]), .Z(n16035) );
  COND1XL U15332 ( .A(n17076), .B(n12997), .C(n16035), .Z(n10515) );
  CANR2X1 U15333 ( .A(n12997), .B(poly12_shifted[22]), .C(n18234), .D(
        Poly12[117]), .Z(n16036) );
  COND1XL U15334 ( .A(n16779), .B(n12997), .C(n16036), .Z(n10526) );
  CANR2X1 U15335 ( .A(n12997), .B(poly12_shifted[16]), .C(n17390), .D(
        Poly12[111]), .Z(n16037) );
  COND1XL U15336 ( .A(n17751), .B(n12997), .C(n16037), .Z(n10532) );
  CANR2X1 U15337 ( .A(n12997), .B(Poly12[20]), .C(n17063), .D(
        poly12_shifted[20]), .Z(n16038) );
  COND1XL U15338 ( .A(n17707), .B(n12997), .C(n16038), .Z(n10512) );
  CANR2X1 U15339 ( .A(n12997), .B(Poly12[30]), .C(n17178), .D(
        poly12_shifted[30]), .Z(n16039) );
  COND1XL U15340 ( .A(n13418), .B(n12997), .C(n16039), .Z(n10502) );
  CANR2X1 U15341 ( .A(n12997), .B(Poly12[22]), .C(n17453), .D(
        poly12_shifted[22]), .Z(n16040) );
  COND1XL U15342 ( .A(n17001), .B(n12997), .C(n16040), .Z(n10510) );
  CANR2X1 U15343 ( .A(n12997), .B(Poly12[28]), .C(n17504), .D(
        poly12_shifted[28]), .Z(n16041) );
  COND1XL U15344 ( .A(n11978), .B(n12997), .C(n16041), .Z(n10504) );
  CANR2X1 U15345 ( .A(n12997), .B(Poly12[27]), .C(n17401), .D(
        poly12_shifted[27]), .Z(n16042) );
  COND1XL U15346 ( .A(n17741), .B(n12997), .C(n16042), .Z(n10505) );
  CANR2X1 U15347 ( .A(n15737), .B(poly3_shifted[42]), .C(n17144), .D(
        poly3_shifted[28]), .Z(n16043) );
  COND1XL U15348 ( .A(n11978), .B(n15737), .C(n16043), .Z(n8912) );
  CANR2X1 U15349 ( .A(n15737), .B(poly3_shifted[22]), .C(n17144), .D(Poly3[78]), .Z(n16044) );
  COND1XL U15350 ( .A(n17163), .B(n15737), .C(n16044), .Z(n8932) );
  CANR2X1 U15351 ( .A(n15737), .B(poly3_shifted[20]), .C(n17144), .D(Poly3[76]), .Z(n16045) );
  COND1XL U15352 ( .A(n16779), .B(n15737), .C(n16045), .Z(n8934) );
  CANR2X1 U15353 ( .A(n15737), .B(poly3_shifted[24]), .C(n17156), .D(Poly3[80]), .Z(n16046) );
  COND1XL U15354 ( .A(n12014), .B(n15737), .C(n16046), .Z(n8930) );
  CANR2X1 U15355 ( .A(n15737), .B(poly3_shifted[14]), .C(n17523), .D(Poly3[70]), .Z(n16047) );
  COND1XL U15356 ( .A(n12011), .B(n15737), .C(n16047), .Z(n8940) );
  CANR2X1 U15357 ( .A(n15737), .B(poly3_shifted[27]), .C(n17144), .D(Poly3[83]), .Z(n16048) );
  COND1XL U15358 ( .A(n17065), .B(n15737), .C(n16048), .Z(n8927) );
  CANR2X1 U15359 ( .A(n15737), .B(poly3_shifted[17]), .C(n17158), .D(Poly3[73]), .Z(n16049) );
  COND1XL U15360 ( .A(n13275), .B(n15737), .C(n16049), .Z(n8937) );
  CANR2X1 U15361 ( .A(n15737), .B(poly3_shifted[31]), .C(n17158), .D(
        poly3_shifted[17]), .Z(n16050) );
  COND1XL U15362 ( .A(n17173), .B(n15737), .C(n16050), .Z(n8923) );
  CANR2X1 U15363 ( .A(n15737), .B(poly3_shifted[44]), .C(n17356), .D(
        poly3_shifted[30]), .Z(n16051) );
  COND1XL U15364 ( .A(n17004), .B(n15737), .C(n16051), .Z(n8910) );
  CANR2X1 U15365 ( .A(n15737), .B(poly3_shifted[38]), .C(n17156), .D(
        poly3_shifted[24]), .Z(n16052) );
  COND1XL U15366 ( .A(n17721), .B(n15737), .C(n16052), .Z(n8916) );
  CANR2X1 U15367 ( .A(n15737), .B(poly3_shifted[16]), .C(n17356), .D(Poly3[72]), .Z(n16053) );
  COND1XL U15368 ( .A(n16303), .B(n15737), .C(n16053), .Z(n8938) );
  CAN2XL U15369 ( .A(n18017), .B(poly8_shifted[57]), .Z(n16054) );
  CANR1XL U15370 ( .A(poly8_shifted[71]), .B(n12287), .C(n16054), .Z(n16055)
         );
  COND1XL U15371 ( .A(n17200), .B(n12287), .C(n16055), .Z(n11344) );
  CANR2X1 U15372 ( .A(n13129), .B(Poly14[177]), .C(n17560), .D(
        poly14_shifted[177]), .Z(n16056) );
  COND1XL U15373 ( .A(n17173), .B(n13129), .C(n16056), .Z(n10228) );
  CANR2X1 U15374 ( .A(n12202), .B(Poly14[206]), .C(n17105), .D(
        poly14_shifted[206]), .Z(n16057) );
  COND1XL U15375 ( .A(n12764), .B(n12202), .C(n16057), .Z(n10199) );
  CANR2X1 U15376 ( .A(n12008), .B(poly14_shifted[158]), .C(n16644), .D(
        poly14_shifted[142]), .Z(n16058) );
  COND1XL U15377 ( .A(n12764), .B(n12008), .C(n16058), .Z(n10263) );
  CANR2X1 U15378 ( .A(n17955), .B(poly9_shifted[89]), .C(n16312), .D(
        poly9_shifted[78]), .Z(n16059) );
  COND1XL U15379 ( .A(n12764), .B(n17955), .C(n16059), .Z(n11227) );
  CEOXL U15380 ( .A(Poly6[47]), .B(Poly6[36]), .Z(n16060) );
  CMXI2X1 U15381 ( .A0(n16957), .A1(n16959), .S(n16060), .Z(n16061) );
  CANR1XL U15382 ( .A(Poly6[46]), .B(n16063), .C(n16061), .Z(n16062) );
  COND1XL U15383 ( .A(n12764), .B(n16063), .C(n16062), .Z(n9647) );
  CANR2X1 U15384 ( .A(n13129), .B(Poly14[174]), .C(n16435), .D(
        poly14_shifted[174]), .Z(n16064) );
  COND1XL U15385 ( .A(n12764), .B(n13129), .C(n16064), .Z(n10231) );
  CANR2X1 U15386 ( .A(n17430), .B(Poly13[526]), .C(n17538), .D(
        poly13_shifted[526]), .Z(n16065) );
  COND1XL U15387 ( .A(n12764), .B(n17430), .C(n16065), .Z(n10534) );
  CANR2X1 U15388 ( .A(n18198), .B(poly1_shifted[313]), .C(n17198), .D(
        poly1_shifted[302]), .Z(n16066) );
  COND1XL U15389 ( .A(n12764), .B(n18198), .C(n16066), .Z(n9055) );
  CENX1 U15390 ( .A(Poly4[59]), .B(Poly4[29]), .Z(n16067) );
  CENX1 U15391 ( .A(n16068), .B(n16067), .Z(n16069) );
  CNR2XL U15392 ( .A(n16069), .B(n17959), .Z(n16070) );
  CANR1XL U15393 ( .A(Poly4[46]), .B(n12153), .C(n16070), .Z(n16071) );
  COND1XL U15394 ( .A(n12764), .B(n12153), .C(n16071), .Z(n8810) );
  CANR2X1 U15395 ( .A(n12185), .B(poly11_shifted[29]), .C(n17552), .D(
        Poly11[85]), .Z(n16072) );
  COND1XL U15396 ( .A(n12764), .B(n12185), .C(n16072), .Z(n11175) );
  CANR2X1 U15397 ( .A(n12009), .B(poly14_shifted[126]), .C(n16644), .D(
        poly14_shifted[110]), .Z(n16073) );
  COND1XL U15398 ( .A(n12764), .B(n12009), .C(n16073), .Z(n10295) );
  CANR2X1 U15399 ( .A(n12262), .B(Poly9[110]), .C(n17545), .D(
        poly9_shifted[110]), .Z(n16074) );
  COND1XL U15400 ( .A(n12764), .B(n12262), .C(n16074), .Z(n11195) );
  CANR2X1 U15401 ( .A(n15737), .B(poly3_shifted[28]), .C(n17375), .D(
        poly3_shifted[14]), .Z(n16075) );
  COND1XL U15402 ( .A(n12764), .B(n15737), .C(n16075), .Z(n8926) );
  CANR2X1 U15403 ( .A(n13351), .B(poly9_shifted[57]), .C(poly9_shifted[46]), 
        .D(n17755), .Z(n16076) );
  COND1XL U15404 ( .A(n12764), .B(n13351), .C(n16076), .Z(n11259) );
  CANR2X1 U15405 ( .A(n12997), .B(poly12_shifted[30]), .C(n17965), .D(
        Poly12[125]), .Z(n16077) );
  COND1XL U15406 ( .A(n12764), .B(n12997), .C(n16077), .Z(n10518) );
  CANR2X1 U15407 ( .A(n17376), .B(Poly15[57]), .C(n17352), .D(
        poly15_shifted[57]), .Z(n16078) );
  COND1XL U15408 ( .A(n17123), .B(n17376), .C(n16078), .Z(n9580) );
  CIVXL U15409 ( .A(poly0_shifted[117]), .Z(n16080) );
  CANR2X1 U15410 ( .A(n18053), .B(n16274), .C(n17352), .D(poly0_shifted[99]), 
        .Z(n16079) );
  COND1XL U15411 ( .A(n16080), .B(n16276), .C(n16079), .Z(n9478) );
  CIVXL U15412 ( .A(Poly0[115]), .Z(n16082) );
  CANR2XL U15413 ( .A(n18176), .B(n16274), .C(n17352), .D(poly0_shifted[115]), 
        .Z(n16081) );
  COND1XL U15414 ( .A(n16082), .B(n16276), .C(n16081), .Z(n9462) );
  CIVXL U15415 ( .A(poly0_shifted[120]), .Z(n16084) );
  CANR2X1 U15416 ( .A(n18116), .B(n16274), .C(n17352), .D(poly0_shifted[102]), 
        .Z(n16083) );
  COND1XL U15417 ( .A(n16084), .B(n16276), .C(n16083), .Z(n9475) );
  CIVX1 U15418 ( .A(Poly0[117]), .Z(n16086) );
  CANR2XL U15419 ( .A(n18241), .B(n16274), .C(n17352), .D(poly0_shifted[117]), 
        .Z(n16085) );
  COND1XL U15420 ( .A(n16086), .B(n16276), .C(n16085), .Z(n9460) );
  CIVXL U15421 ( .A(Poly0[120]), .Z(n16088) );
  CANR2X1 U15422 ( .A(n13994), .B(n16274), .C(n17352), .D(poly0_shifted[120]), 
        .Z(n16087) );
  COND1XL U15423 ( .A(n16088), .B(n16276), .C(n16087), .Z(n9457) );
  CANR2X1 U15424 ( .A(n12008), .B(poly14_shifted[172]), .C(n17642), .D(
        poly14_shifted[156]), .Z(n16089) );
  COND1XL U15425 ( .A(n11978), .B(n12008), .C(n16089), .Z(n10249) );
  CANR2X1 U15426 ( .A(n12009), .B(poly14_shifted[140]), .C(n17965), .D(
        poly14_shifted[124]), .Z(n16090) );
  COND1XL U15427 ( .A(n11978), .B(n12009), .C(n16090), .Z(n10281) );
  CAOR1X1 U15428 ( .A(n16091), .B(n16094), .C(n18219), .Z(n16092) );
  CMXI2X1 U15429 ( .A0(n16092), .A1(Poly10[13]), .S(n17962), .Z(n16093) );
  COND11XL U15430 ( .A(Poly10[39]), .B(n17495), .C(n16094), .D(n16093), .Z(
        n11090) );
  CANR2X1 U15431 ( .A(n12977), .B(poly7_shifted[178]), .C(n17620), .D(
        poly7_shifted[166]), .Z(n16095) );
  COND1XL U15432 ( .A(n17757), .B(n12977), .C(n16095), .Z(n9938) );
  CANR2X1 U15433 ( .A(n16425), .B(poly1_shifted[109]), .C(n17334), .D(
        poly1_shifted[98]), .Z(n16096) );
  COND1XL U15434 ( .A(n16775), .B(n16425), .C(n16096), .Z(n9259) );
  CANR2X1 U15435 ( .A(n16425), .B(poly1_shifted[137]), .C(n18234), .D(
        poly1_shifted[126]), .Z(n16097) );
  COND1XL U15436 ( .A(n17004), .B(n16425), .C(n16097), .Z(n9231) );
  CANR2X1 U15437 ( .A(n16425), .B(poly1_shifted[117]), .C(n18047), .D(
        poly1_shifted[106]), .Z(n16098) );
  COND1XL U15438 ( .A(n12014), .B(n16425), .C(n16098), .Z(n9251) );
  CANR2X1 U15439 ( .A(n16425), .B(poly1_shifted[131]), .C(n17343), .D(
        poly1_shifted[120]), .Z(n16099) );
  COND1XL U15440 ( .A(n17721), .B(n16425), .C(n16099), .Z(n9237) );
  CANR2X1 U15441 ( .A(n16425), .B(poly1_shifted[122]), .C(n17705), .D(
        poly1_shifted[111]), .Z(n16100) );
  COND1XL U15442 ( .A(n17196), .B(n16425), .C(n16100), .Z(n9246) );
  CANR2X1 U15443 ( .A(n16425), .B(poly1_shifted[120]), .C(n17655), .D(
        poly1_shifted[109]), .Z(n16101) );
  COND1XL U15444 ( .A(n17090), .B(n16425), .C(n16101), .Z(n9248) );
  CANR2X1 U15445 ( .A(n16425), .B(poly1_shifted[134]), .C(n18234), .D(
        poly1_shifted[123]), .Z(n16102) );
  COND1XL U15446 ( .A(n17741), .B(n16425), .C(n16102), .Z(n9234) );
  CANR2X1 U15447 ( .A(n16425), .B(poly1_shifted[112]), .C(n17640), .D(
        poly1_shifted[101]), .Z(n16103) );
  COND1XL U15448 ( .A(n11993), .B(n16425), .C(n16103), .Z(n9256) );
  CANR2X1 U15449 ( .A(n17974), .B(poly13_shifted[138]), .C(n17755), .D(
        poly13_shifted[124]), .Z(n16104) );
  COND1XL U15450 ( .A(n11978), .B(n17974), .C(n16104), .Z(n10936) );
  CANR2X1 U15451 ( .A(n17987), .B(poly13_shifted[430]), .C(n18047), .D(
        poly13_shifted[416]), .Z(n16105) );
  COND1XL U15452 ( .A(n12011), .B(n17987), .C(n16105), .Z(n10644) );
  CANR2X1 U15453 ( .A(n17987), .B(poly13_shifted[455]), .C(n17552), .D(
        poly13_shifted[441]), .Z(n16106) );
  COND1XL U15454 ( .A(n17200), .B(n17987), .C(n16106), .Z(n10619) );
  CANR2X1 U15455 ( .A(n17987), .B(poly13_shifted[444]), .C(n18017), .D(
        poly13_shifted[430]), .Z(n16107) );
  COND1XL U15456 ( .A(n12764), .B(n17987), .C(n16107), .Z(n10630) );
  CANR2X1 U15457 ( .A(n17982), .B(poly13_shifted[393]), .C(n16427), .D(
        poly13_shifted[379]), .Z(n16108) );
  COND1XL U15458 ( .A(n17741), .B(n17982), .C(n16108), .Z(n10681) );
  CANR2X1 U15459 ( .A(n17987), .B(poly13_shifted[431]), .C(n17458), .D(
        poly13_shifted[417]), .Z(n16109) );
  COND1XL U15460 ( .A(n16950), .B(n17987), .C(n16109), .Z(n10643) );
  CANR2X1 U15461 ( .A(n17982), .B(poly13_shifted[375]), .C(n17755), .D(
        poly13_shifted[361]), .Z(n16110) );
  COND1XL U15462 ( .A(n17208), .B(n17982), .C(n16110), .Z(n10699) );
  CANR2X1 U15463 ( .A(n17982), .B(poly13_shifted[391]), .C(n17466), .D(
        poly13_shifted[377]), .Z(n16111) );
  COND1XL U15464 ( .A(n17200), .B(n17982), .C(n16111), .Z(n10683) );
  CANR2X1 U15465 ( .A(n17982), .B(poly13_shifted[376]), .C(n17755), .D(
        poly13_shifted[362]), .Z(n16112) );
  COND1XL U15466 ( .A(n12014), .B(n17982), .C(n16112), .Z(n10698) );
  CANR2X1 U15467 ( .A(n17974), .B(poly13_shifted[111]), .C(n17348), .D(
        poly13_shifted[97]), .Z(n16113) );
  COND1XL U15468 ( .A(n16950), .B(n17974), .C(n16113), .Z(n10963) );
  CANR2X1 U15469 ( .A(n17982), .B(poly13_shifted[394]), .C(n17705), .D(
        poly13_shifted[380]), .Z(n16114) );
  COND1XL U15470 ( .A(n11978), .B(n17982), .C(n16114), .Z(n10680) );
  CANR2X1 U15471 ( .A(n17974), .B(poly13_shifted[137]), .C(n16787), .D(
        poly13_shifted[123]), .Z(n16115) );
  COND1XL U15472 ( .A(n17741), .B(n17974), .C(n16115), .Z(n10937) );
  CANR2X1 U15473 ( .A(n17987), .B(poly13_shifted[442]), .C(n17383), .D(
        poly13_shifted[428]), .Z(n16116) );
  COND1XL U15474 ( .A(n17087), .B(n17987), .C(n16116), .Z(n10632) );
  CANR2X1 U15475 ( .A(n17982), .B(poly13_shifted[380]), .C(n17121), .D(
        poly13_shifted[366]), .Z(n16117) );
  COND1XL U15476 ( .A(n17699), .B(n17982), .C(n16117), .Z(n10694) );
  CANR2X1 U15477 ( .A(n17987), .B(poly13_shifted[443]), .C(n17755), .D(
        poly13_shifted[429]), .Z(n16118) );
  COND1XL U15478 ( .A(n17090), .B(n17987), .C(n16118), .Z(n10631) );
  CANR2X1 U15479 ( .A(n17974), .B(poly13_shifted[122]), .C(n17280), .D(
        poly13_shifted[108]), .Z(n16119) );
  COND1XL U15480 ( .A(n17087), .B(n17974), .C(n16119), .Z(n10952) );
  CANR2X1 U15481 ( .A(n17974), .B(poly13_shifted[125]), .C(n17538), .D(
        poly13_shifted[111]), .Z(n16120) );
  COND1XL U15482 ( .A(n17196), .B(n17974), .C(n16120), .Z(n10949) );
  CANR2X1 U15483 ( .A(n17974), .B(poly13_shifted[139]), .C(n17545), .D(
        poly13_shifted[125]), .Z(n16121) );
  COND1XL U15484 ( .A(n17185), .B(n17974), .C(n16121), .Z(n10935) );
  CANR2X1 U15485 ( .A(n17982), .B(poly13_shifted[381]), .C(n17634), .D(
        poly13_shifted[367]), .Z(n16122) );
  COND1XL U15486 ( .A(n17196), .B(n17982), .C(n16122), .Z(n10693) );
  CANR2X1 U15487 ( .A(n12009), .B(poly14_shifted[137]), .C(n16695), .D(
        poly14_shifted[121]), .Z(n16123) );
  COND1XL U15488 ( .A(n17123), .B(n12009), .C(n16123), .Z(n10284) );
  CAN2XL U15489 ( .A(n18017), .B(poly12_shifted[57]), .Z(n16124) );
  CANR1XL U15490 ( .A(Poly12[57]), .B(n12598), .C(n16124), .Z(n16125) );
  COND1XL U15491 ( .A(n17123), .B(n12598), .C(n16125), .Z(n10475) );
  CANR2X1 U15492 ( .A(n12932), .B(poly14_shifted[297]), .C(n17545), .D(
        poly14_shifted[281]), .Z(n16126) );
  COND1XL U15493 ( .A(n17123), .B(n12932), .C(n16126), .Z(n10124) );
  CANR2X1 U15494 ( .A(n18018), .B(poly7_shifted[14]), .C(n17209), .D(
        Poly7[401]), .Z(n16127) );
  COND1XL U15495 ( .A(n16303), .B(n18018), .C(n16127), .Z(n10102) );
  CANR2X1 U15496 ( .A(n17273), .B(poly7_shifted[229]), .C(n16695), .D(
        poly7_shifted[217]), .Z(n16128) );
  COND1XL U15497 ( .A(n17200), .B(n17273), .C(n16128), .Z(n9887) );
  CANR2X1 U15498 ( .A(n17273), .B(poly7_shifted[231]), .C(n17466), .D(
        poly7_shifted[219]), .Z(n16129) );
  COND1XL U15499 ( .A(n17741), .B(n17273), .C(n16129), .Z(n9885) );
  CANR2X1 U15500 ( .A(n17273), .B(poly7_shifted[235]), .C(n17705), .D(
        poly7_shifted[223]), .Z(n16130) );
  COND1XL U15501 ( .A(n17188), .B(n17273), .C(n16130), .Z(n9881) );
  CANR2X1 U15502 ( .A(n12009), .B(poly14_shifted[113]), .C(n17488), .D(
        poly14_shifted[97]), .Z(n16131) );
  COND1XL U15503 ( .A(n16950), .B(n12009), .C(n16131), .Z(n10308) );
  CANR2X1 U15504 ( .A(n12008), .B(poly14_shifted[145]), .C(n18234), .D(
        poly14_shifted[129]), .Z(n16132) );
  COND1XL U15505 ( .A(n16950), .B(n12008), .C(n16132), .Z(n10276) );
  CANR2X1 U15506 ( .A(n13129), .B(poly14_shifted[177]), .C(n17552), .D(
        poly14_shifted[161]), .Z(n16133) );
  COND1XL U15507 ( .A(n16950), .B(n13129), .C(n16133), .Z(n10244) );
  CANR2XL U15508 ( .A(n12932), .B(poly14_shifted[273]), .C(n17998), .D(
        poly14_shifted[257]), .Z(n16134) );
  COND1XL U15509 ( .A(n16950), .B(n12932), .C(n16134), .Z(n10148) );
  CEOX1 U15510 ( .A(n16135), .B(n18238), .Z(n16136) );
  CEOX1 U15511 ( .A(n16136), .B(dataselector[49]), .Z(n16137) );
  CANR2X1 U15512 ( .A(n16350), .B(dataselector[56]), .C(n16137), .D(n18017), 
        .Z(n16138) );
  COND1XL U15513 ( .A(n16139), .B(n17721), .C(n16138), .Z(n8739) );
  CANR2X1 U15514 ( .A(n18018), .B(poly7_shifted[27]), .C(n17383), .D(
        poly7_shifted[15]), .Z(n16140) );
  COND1XL U15515 ( .A(n17196), .B(n18018), .C(n16140), .Z(n10089) );
  CANR2X1 U15516 ( .A(n18018), .B(poly7_shifted[29]), .C(n17209), .D(
        poly7_shifted[17]), .Z(n16141) );
  COND1XL U15517 ( .A(n17173), .B(n18018), .C(n16141), .Z(n10087) );
  CANR2X1 U15518 ( .A(n18018), .B(Poly7[27]), .C(n17383), .D(poly7_shifted[27]), .Z(n16142) );
  COND1XL U15519 ( .A(n17741), .B(n18018), .C(n16142), .Z(n10077) );
  CANR2X1 U15520 ( .A(n17974), .B(poly13_shifted[117]), .C(n17488), .D(
        poly13_shifted[103]), .Z(n16143) );
  COND1XL U15521 ( .A(n16939), .B(n17974), .C(n16143), .Z(n10957) );
  CANR2X1 U15522 ( .A(n17987), .B(poly13_shifted[460]), .C(n17755), .D(
        poly13_shifted[446]), .Z(n16144) );
  COND1XL U15523 ( .A(n13418), .B(n17987), .C(n16144), .Z(n10614) );
  CANR2X1 U15524 ( .A(n17987), .B(poly13_shifted[437]), .C(poly13_shifted[423]), .D(n17755), .Z(n16145) );
  COND1XL U15525 ( .A(n17718), .B(n17987), .C(n16145), .Z(n10637) );
  CANR2X1 U15526 ( .A(n17974), .B(poly13_shifted[119]), .C(n17642), .D(
        poly13_shifted[105]), .Z(n16146) );
  COND1XL U15527 ( .A(n17208), .B(n17974), .C(n16146), .Z(n10955) );
  CANR2X1 U15528 ( .A(n17974), .B(poly13_shifted[116]), .C(n17620), .D(
        poly13_shifted[102]), .Z(n16147) );
  COND1XL U15529 ( .A(n16779), .B(n17974), .C(n16147), .Z(n10958) );
  CANR2X1 U15530 ( .A(n17982), .B(poly13_shifted[386]), .C(n17640), .D(
        poly13_shifted[372]), .Z(n16148) );
  COND1XL U15531 ( .A(n17707), .B(n17982), .C(n16148), .Z(n10688) );
  CANR2X1 U15532 ( .A(n17982), .B(poly13_shifted[397]), .C(n17238), .D(
        poly13_shifted[383]), .Z(n16149) );
  COND1XL U15533 ( .A(n17188), .B(n17982), .C(n16149), .Z(n10677) );
  CANR2X1 U15534 ( .A(n17974), .B(poly13_shifted[112]), .C(n16435), .D(
        poly13_shifted[98]), .Z(n16150) );
  COND1XL U15535 ( .A(n16775), .B(n17974), .C(n16150), .Z(n10962) );
  CANR2X1 U15536 ( .A(n17974), .B(poly13_shifted[140]), .C(n17640), .D(
        poly13_shifted[126]), .Z(n16151) );
  COND1XL U15537 ( .A(n13418), .B(n17974), .C(n16151), .Z(n10934) );
  CANR2X1 U15538 ( .A(n17974), .B(poly13_shifted[126]), .C(n17295), .D(
        poly13_shifted[112]), .Z(n16152) );
  COND1XL U15539 ( .A(n17062), .B(n17974), .C(n16152), .Z(n10948) );
  CANR2X1 U15540 ( .A(n17982), .B(poly13_shifted[369]), .C(n17072), .D(
        poly13_shifted[355]), .Z(n16153) );
  COND1XL U15541 ( .A(n13275), .B(n17982), .C(n16153), .Z(n10705) );
  CANR2X1 U15542 ( .A(n17982), .B(poly13_shifted[388]), .C(n17965), .D(
        poly13_shifted[374]), .Z(n16154) );
  COND1XL U15543 ( .A(n17001), .B(n17982), .C(n16154), .Z(n10686) );
  CANR2X1 U15544 ( .A(n17982), .B(poly13_shifted[383]), .C(n17449), .D(
        poly13_shifted[369]), .Z(n16155) );
  COND1XL U15545 ( .A(n17173), .B(n17982), .C(n16155), .Z(n10691) );
  CANR2X1 U15546 ( .A(n17974), .B(poly13_shifted[132]), .C(n17298), .D(
        poly13_shifted[118]), .Z(n16156) );
  COND1XL U15547 ( .A(n17001), .B(n17974), .C(n16156), .Z(n10942) );
  CANR2X1 U15548 ( .A(n17982), .B(poly13_shifted[378]), .C(n17620), .D(
        poly13_shifted[364]), .Z(n16157) );
  COND1XL U15549 ( .A(n17087), .B(n17982), .C(n16157), .Z(n10696) );
  CANR2X1 U15550 ( .A(n17974), .B(poly13_shifted[131]), .C(n17401), .D(
        poly13_shifted[117]), .Z(n16158) );
  COND1XL U15551 ( .A(n12006), .B(n17974), .C(n16158), .Z(n10943) );
  CANR2X1 U15552 ( .A(n17982), .B(poly13_shifted[395]), .C(n17620), .D(
        poly13_shifted[381]), .Z(n16159) );
  COND1XL U15553 ( .A(n17185), .B(n17982), .C(n16159), .Z(n10679) );
  CANR2X1 U15554 ( .A(n17982), .B(poly13_shifted[377]), .C(n17466), .D(
        poly13_shifted[363]), .Z(n16160) );
  COND1XL U15555 ( .A(n16605), .B(n17982), .C(n16160), .Z(n10697) );
  CANR2X1 U15556 ( .A(n17987), .B(poly13_shifted[458]), .C(n17508), .D(
        poly13_shifted[444]), .Z(n16161) );
  COND1XL U15557 ( .A(n11978), .B(n17987), .C(n16161), .Z(n10616) );
  CANR2X1 U15558 ( .A(n17982), .B(poly13_shifted[396]), .C(n16583), .D(
        poly13_shifted[382]), .Z(n16162) );
  COND1XL U15559 ( .A(n13418), .B(n17982), .C(n16162), .Z(n10678) );
  CANR2X1 U15560 ( .A(n17987), .B(poly13_shifted[440]), .C(n17508), .D(
        poly13_shifted[426]), .Z(n16163) );
  COND1XL U15561 ( .A(n12014), .B(n17987), .C(n16163), .Z(n10634) );
  CANR2X1 U15562 ( .A(n17982), .B(poly13_shifted[367]), .C(n16488), .D(
        poly13_shifted[353]), .Z(n16164) );
  COND1XL U15563 ( .A(n17697), .B(n17982), .C(n16164), .Z(n10707) );
  CANR2X1 U15564 ( .A(n17982), .B(poly13_shifted[382]), .C(n17158), .D(
        poly13_shifted[368]), .Z(n16165) );
  COND1XL U15565 ( .A(n17062), .B(n17982), .C(n16165), .Z(n10692) );
  CANR2X1 U15566 ( .A(n17987), .B(poly13_shifted[454]), .C(n17390), .D(
        poly13_shifted[440]), .Z(n16166) );
  COND1XL U15567 ( .A(n17721), .B(n17987), .C(n16166), .Z(n10620) );
  CANR2X1 U15568 ( .A(n17987), .B(poly13_shifted[438]), .C(n17755), .D(
        poly13_shifted[424]), .Z(n16167) );
  COND1XL U15569 ( .A(n17163), .B(n17987), .C(n16167), .Z(n10636) );
  CANR2X1 U15570 ( .A(n17974), .B(poly13_shifted[127]), .C(n17348), .D(
        poly13_shifted[113]), .Z(n16168) );
  COND1XL U15571 ( .A(n17076), .B(n17974), .C(n16168), .Z(n10947) );
  CANR2X1 U15572 ( .A(n17974), .B(poly13_shifted[110]), .C(n17348), .D(
        poly13_shifted[96]), .Z(n16169) );
  COND1XL U15573 ( .A(n17751), .B(n17974), .C(n16169), .Z(n10964) );
  CANR2X1 U15574 ( .A(n17982), .B(poly13_shifted[368]), .C(n17398), .D(
        poly13_shifted[354]), .Z(n16170) );
  COND1XL U15575 ( .A(n16775), .B(n17982), .C(n16170), .Z(n10706) );
  CANR2X1 U15576 ( .A(n17974), .B(poly13_shifted[113]), .C(n18234), .D(
        poly13_shifted[99]), .Z(n16171) );
  COND1XL U15577 ( .A(n13275), .B(n17974), .C(n16171), .Z(n10961) );
  CANR2X1 U15578 ( .A(n17987), .B(poly13_shifted[432]), .C(n16583), .D(
        poly13_shifted[418]), .Z(n16172) );
  COND1XL U15579 ( .A(n16775), .B(n17987), .C(n16172), .Z(n10642) );
  CANR2X1 U15580 ( .A(n17974), .B(poly13_shifted[121]), .C(n17755), .D(
        poly13_shifted[107]), .Z(n16173) );
  COND1XL U15581 ( .A(n16994), .B(n17974), .C(n16173), .Z(n10953) );
  CANR2X1 U15582 ( .A(n17987), .B(poly13_shifted[445]), .C(n17453), .D(
        poly13_shifted[431]), .Z(n16174) );
  COND1XL U15583 ( .A(n17196), .B(n17987), .C(n16174), .Z(n10629) );
  CANR2X1 U15584 ( .A(n17987), .B(poly13_shifted[441]), .C(n18234), .D(
        poly13_shifted[427]), .Z(n16175) );
  COND1XL U15585 ( .A(n16994), .B(n17987), .C(n16175), .Z(n10633) );
  CANR2X1 U15586 ( .A(n17974), .B(poly13_shifted[123]), .C(n17705), .D(
        poly13_shifted[109]), .Z(n16176) );
  COND1XL U15587 ( .A(n17065), .B(n17974), .C(n16176), .Z(n10951) );
  CANR2X1 U15588 ( .A(n17987), .B(poly13_shifted[450]), .C(n16583), .D(
        poly13_shifted[436]), .Z(n16177) );
  COND1XL U15589 ( .A(n17707), .B(n17987), .C(n16177), .Z(n10624) );
  CANR2X1 U15590 ( .A(n17974), .B(poly13_shifted[134]), .C(n17755), .D(
        poly13_shifted[120]), .Z(n16178) );
  COND1XL U15591 ( .A(n16179), .B(n17974), .C(n16178), .Z(n10940) );
  CANR2XL U15592 ( .A(n17667), .B(poly13_shifted[207]), .C(n17285), .D(
        poly13_shifted[193]), .Z(n16180) );
  COND1XL U15593 ( .A(n16950), .B(n17667), .C(n16180), .Z(n10867) );
  CANR2XL U15594 ( .A(n17667), .B(poly13_shifted[221]), .C(n17285), .D(
        poly13_shifted[207]), .Z(n16181) );
  COND1XL U15595 ( .A(n17196), .B(n17667), .C(n16181), .Z(n10853) );
  CANR2X1 U15596 ( .A(n13014), .B(poly13_shifted[199]), .C(n17449), .D(
        poly13_shifted[185]), .Z(n16182) );
  COND1XL U15597 ( .A(n17200), .B(n13014), .C(n16182), .Z(n10875) );
  CANR2X1 U15598 ( .A(n13014), .B(poly13_shifted[204]), .C(n17285), .D(
        poly13_shifted[190]), .Z(n16183) );
  COND1XL U15599 ( .A(n13418), .B(n13014), .C(n16183), .Z(n10870) );
  CANR2X1 U15600 ( .A(n13014), .B(poly13_shifted[203]), .C(n17094), .D(
        poly13_shifted[189]), .Z(n16184) );
  COND1XL U15601 ( .A(n17185), .B(n13014), .C(n16184), .Z(n10871) );
  CEOXL U15602 ( .A(Poly13[519]), .B(Poly13[160]), .Z(n16185) );
  CANR2X1 U15603 ( .A(n13014), .B(poly13_shifted[188]), .C(n17998), .D(n16185), 
        .Z(n16186) );
  COND1XL U15604 ( .A(n12764), .B(n13014), .C(n16186), .Z(n10886) );
  CEOXL U15605 ( .A(Poly13[518]), .B(Poly13[159]), .Z(n16187) );
  CANR2X1 U15606 ( .A(n13014), .B(poly13_shifted[187]), .C(n17362), .D(n16187), 
        .Z(n16188) );
  COND1XL U15607 ( .A(n17065), .B(n13014), .C(n16188), .Z(n10887) );
  CANR2X1 U15608 ( .A(n13014), .B(Poly13[160]), .C(n17508), .D(
        poly13_shifted[160]), .Z(n16189) );
  COND1XL U15609 ( .A(n17751), .B(n13014), .C(n16189), .Z(n10900) );
  CANR2X1 U15610 ( .A(n13014), .B(poly13_shifted[198]), .C(n18234), .D(
        poly13_shifted[184]), .Z(n16190) );
  COND1XL U15611 ( .A(n17721), .B(n13014), .C(n16190), .Z(n10876) );
  CANR2X1 U15612 ( .A(n13014), .B(poly13_shifted[201]), .C(n16427), .D(
        poly13_shifted[187]), .Z(n16191) );
  COND1XL U15613 ( .A(n17741), .B(n13014), .C(n16191), .Z(n10873) );
  CANR2X1 U15614 ( .A(n17603), .B(poly13_shifted[350]), .C(n17755), .D(
        poly13_shifted[336]), .Z(n16192) );
  COND1XL U15615 ( .A(n17062), .B(n17603), .C(n16192), .Z(n10724) );
  CANR2X1 U15616 ( .A(n18002), .B(poly14_shifted[27]), .C(n16999), .D(
        Poly14[296]), .Z(n16193) );
  COND1XL U15617 ( .A(n16605), .B(n18002), .C(n16193), .Z(n10394) );
  CANR2X1 U15618 ( .A(n18002), .B(poly14_shifted[43]), .C(n16999), .D(
        poly14_shifted[27]), .Z(n16194) );
  COND1XL U15619 ( .A(n17741), .B(n18002), .C(n16194), .Z(n10378) );
  CANR2X1 U15620 ( .A(n13014), .B(Poly13[161]), .C(n17642), .D(
        poly13_shifted[161]), .Z(n16195) );
  COND1XL U15621 ( .A(n16950), .B(n13014), .C(n16195), .Z(n10899) );
  CANR2X1 U15622 ( .A(n13014), .B(Poly13[162]), .C(n17755), .D(
        poly13_shifted[162]), .Z(n16196) );
  COND1XL U15623 ( .A(n16775), .B(n13014), .C(n16196), .Z(n10898) );
  CANR2X1 U15624 ( .A(n13014), .B(poly13_shifted[205]), .C(n17755), .D(
        poly13_shifted[191]), .Z(n16197) );
  COND1XL U15625 ( .A(n17188), .B(n13014), .C(n16197), .Z(n10869) );
  CANR2X1 U15626 ( .A(n13014), .B(Poly13[167]), .C(n18234), .D(
        poly13_shifted[167]), .Z(n16198) );
  COND1XL U15627 ( .A(n16939), .B(n13014), .C(n16198), .Z(n10893) );
  CEOXL U15628 ( .A(Poly14[294]), .B(Poly14[300]), .Z(n16199) );
  CENX1 U15629 ( .A(Poly14[208]), .B(n16199), .Z(n16200) );
  CNR2X1 U15630 ( .A(n16200), .B(n17495), .Z(n16201) );
  CANR1XL U15631 ( .A(poly14_shifted[240]), .B(n16694), .C(n16201), .Z(n16202)
         );
  COND1XL U15632 ( .A(n12011), .B(n16694), .C(n16202), .Z(n10181) );
  CANR2X1 U15633 ( .A(n17273), .B(poly7_shifted[234]), .C(n17535), .D(
        poly7_shifted[222]), .Z(n16203) );
  COND1XL U15634 ( .A(n13418), .B(n17273), .C(n16203), .Z(n9882) );
  CANR2X1 U15635 ( .A(n17273), .B(poly7_shifted[225]), .C(n16488), .D(
        poly7_shifted[213]), .Z(n16204) );
  COND1XL U15636 ( .A(n12006), .B(n17273), .C(n16204), .Z(n9891) );
  CANR2X1 U15637 ( .A(n17273), .B(poly7_shifted[233]), .C(n17533), .D(
        poly7_shifted[221]), .Z(n16205) );
  COND1XL U15638 ( .A(n17185), .B(n17273), .C(n16205), .Z(n9883) );
  CANR2X1 U15639 ( .A(n17525), .B(poly14_shifted[63]), .C(n17552), .D(
        poly14_shifted[47]), .Z(n16206) );
  COND1XL U15640 ( .A(n17196), .B(n17525), .C(n16206), .Z(n10358) );
  CANR2X1 U15641 ( .A(n17525), .B(poly14_shifted[49]), .C(n17504), .D(
        poly14_shifted[33]), .Z(n16207) );
  COND1XL U15642 ( .A(n16950), .B(n17525), .C(n16207), .Z(n10372) );
  CANR2X1 U15643 ( .A(n17525), .B(poly14_shifted[72]), .C(n16787), .D(
        poly14_shifted[56]), .Z(n16208) );
  COND1XL U15644 ( .A(n16179), .B(n17525), .C(n16208), .Z(n10349) );
  CANR2X1 U15645 ( .A(n17525), .B(poly14_shifted[65]), .C(n17998), .D(
        poly14_shifted[49]), .Z(n16209) );
  COND1XL U15646 ( .A(n17076), .B(n17525), .C(n16209), .Z(n10356) );
  CANR2X1 U15647 ( .A(n17525), .B(poly14_shifted[70]), .C(n17714), .D(
        poly14_shifted[54]), .Z(n16210) );
  COND1XL U15648 ( .A(n17001), .B(n17525), .C(n16210), .Z(n10351) );
  CANR2X1 U15649 ( .A(n17525), .B(poly14_shifted[57]), .C(n17362), .D(
        poly14_shifted[41]), .Z(n16211) );
  COND1XL U15650 ( .A(n17208), .B(n17525), .C(n16211), .Z(n10364) );
  CANR2X1 U15651 ( .A(n17525), .B(poly14_shifted[50]), .C(n17523), .D(
        poly14_shifted[34]), .Z(n16212) );
  COND1XL U15652 ( .A(n16303), .B(n17525), .C(n16212), .Z(n10371) );
  CANR2X1 U15653 ( .A(n17525), .B(poly14_shifted[48]), .C(n16307), .D(
        poly14_shifted[32]), .Z(n16213) );
  COND1XL U15654 ( .A(n12011), .B(n17525), .C(n16213), .Z(n10373) );
  CANR2XL U15655 ( .A(n17525), .B(poly14_shifted[58]), .C(n18017), .D(
        poly14_shifted[42]), .Z(n16214) );
  COND1XL U15656 ( .A(n12014), .B(n17525), .C(n16214), .Z(n10363) );
  CANR2X1 U15657 ( .A(n17525), .B(poly14_shifted[73]), .C(n16427), .D(
        poly14_shifted[57]), .Z(n16215) );
  COND1XL U15658 ( .A(n17123), .B(n17525), .C(n16215), .Z(n10348) );
  CANR2X1 U15659 ( .A(n17525), .B(poly14_shifted[77]), .C(n17552), .D(
        poly14_shifted[61]), .Z(n16216) );
  COND1XL U15660 ( .A(n17185), .B(n17525), .C(n16216), .Z(n10344) );
  CANR2X1 U15661 ( .A(n17525), .B(poly14_shifted[62]), .C(n16307), .D(
        poly14_shifted[46]), .Z(n16217) );
  COND1XL U15662 ( .A(n12764), .B(n17525), .C(n16217), .Z(n10359) );
  CANR2X1 U15663 ( .A(n17525), .B(poly14_shifted[76]), .C(n17466), .D(
        poly14_shifted[60]), .Z(n16218) );
  COND1XL U15664 ( .A(n11978), .B(n17525), .C(n16218), .Z(n10345) );
  CANR2X1 U15665 ( .A(n17525), .B(poly14_shifted[64]), .C(n17545), .D(
        poly14_shifted[48]), .Z(n16219) );
  COND1XL U15666 ( .A(n17062), .B(n17525), .C(n16219), .Z(n10357) );
  CANR2X1 U15667 ( .A(n17525), .B(poly14_shifted[79]), .C(n16702), .D(
        poly14_shifted[63]), .Z(n16220) );
  COND1XL U15668 ( .A(n17188), .B(n17525), .C(n16220), .Z(n10342) );
  CANR2X1 U15669 ( .A(n17525), .B(poly14_shifted[51]), .C(n17705), .D(
        poly14_shifted[35]), .Z(n16221) );
  COND1XL U15670 ( .A(n13275), .B(n17525), .C(n16221), .Z(n10370) );
  CANR2X1 U15671 ( .A(n17525), .B(poly14_shifted[61]), .C(n18234), .D(
        poly14_shifted[45]), .Z(n16222) );
  COND1XL U15672 ( .A(n17090), .B(n17525), .C(n16222), .Z(n10360) );
  CANR2X1 U15673 ( .A(n17525), .B(poly14_shifted[78]), .C(n16427), .D(
        poly14_shifted[62]), .Z(n16223) );
  COND1XL U15674 ( .A(n17004), .B(n17525), .C(n16223), .Z(n10343) );
  CANR2X1 U15675 ( .A(n17592), .B(Poly13[271]), .C(n17298), .D(
        poly13_shifted[271]), .Z(n16224) );
  COND1XL U15676 ( .A(n17196), .B(n17592), .C(n16224), .Z(n10789) );
  CANR2X1 U15677 ( .A(n17592), .B(poly13_shifted[272]), .C(n17298), .D(
        poly13_shifted[258]), .Z(n16225) );
  COND1XL U15678 ( .A(n16775), .B(n17592), .C(n16225), .Z(n10802) );
  CANR2X1 U15679 ( .A(n17592), .B(poly13_shifted[280]), .C(n18234), .D(
        poly13_shifted[266]), .Z(n16226) );
  COND1XL U15680 ( .A(n12014), .B(n17592), .C(n16226), .Z(n10794) );
  CANR2X1 U15681 ( .A(n17592), .B(poly13_shifted[271]), .C(n17298), .D(
        poly13_shifted[257]), .Z(n16227) );
  COND1XL U15682 ( .A(n16950), .B(n17592), .C(n16227), .Z(n10803) );
  CEOXL U15683 ( .A(Poly13[517]), .B(Poly13[272]), .Z(n16228) );
  CANR2X1 U15684 ( .A(n17592), .B(poly13_shifted[300]), .C(n17298), .D(n16228), 
        .Z(n16229) );
  COND1XL U15685 ( .A(n13418), .B(n17592), .C(n16229), .Z(n10774) );
  CANR2X1 U15686 ( .A(n17592), .B(Poly13[269]), .C(n18234), .D(
        poly13_shifted[269]), .Z(n16230) );
  COND1XL U15687 ( .A(n17090), .B(n17592), .C(n16230), .Z(n10791) );
  CEOXL U15688 ( .A(Poly13[516]), .B(Poly13[271]), .Z(n16231) );
  CANR2X1 U15689 ( .A(n17592), .B(poly13_shifted[299]), .C(n17298), .D(n16231), 
        .Z(n16232) );
  COND1XL U15690 ( .A(n17185), .B(n17592), .C(n16232), .Z(n10775) );
  CANR2X1 U15691 ( .A(n17592), .B(Poly13[272]), .C(n17298), .D(
        poly13_shifted[272]), .Z(n16233) );
  COND1XL U15692 ( .A(n17062), .B(n17592), .C(n16233), .Z(n10788) );
  CANR2X1 U15693 ( .A(n17592), .B(poly13_shifted[270]), .C(n17266), .D(
        poly13_shifted[256]), .Z(n16234) );
  COND1XL U15694 ( .A(n12011), .B(n17592), .C(n16234), .Z(n10804) );
  CANR2X1 U15695 ( .A(n17491), .B(poly13_shifted[524]), .C(n17401), .D(
        poly13_shifted[510]), .Z(n16235) );
  COND1XL U15696 ( .A(n13418), .B(n17491), .C(n16235), .Z(n10550) );
  CANR2X1 U15697 ( .A(n17491), .B(poly13_shifted[505]), .C(n17121), .D(
        poly13_shifted[491]), .Z(n16236) );
  COND1XL U15698 ( .A(n16994), .B(n17491), .C(n16236), .Z(n10569) );
  CANR2X1 U15699 ( .A(n17491), .B(poly13_shifted[495]), .C(n16583), .D(
        poly13_shifted[481]), .Z(n16237) );
  COND1XL U15700 ( .A(n17697), .B(n17491), .C(n16237), .Z(n10579) );
  CANR2X1 U15701 ( .A(n17491), .B(poly13_shifted[516]), .C(n17998), .D(
        poly13_shifted[502]), .Z(n16238) );
  COND1XL U15702 ( .A(n17753), .B(n17491), .C(n16238), .Z(n10558) );
  CANR2X1 U15703 ( .A(n17491), .B(poly13_shifted[506]), .C(n16702), .D(
        poly13_shifted[492]), .Z(n16239) );
  COND1XL U15704 ( .A(n17087), .B(n17491), .C(n16239), .Z(n10568) );
  CANR2X1 U15705 ( .A(n17491), .B(poly13_shifted[523]), .C(n17668), .D(
        poly13_shifted[509]), .Z(n16240) );
  COND1XL U15706 ( .A(n17185), .B(n17491), .C(n16240), .Z(n10551) );
  CANR2X1 U15707 ( .A(n17491), .B(poly13_shifted[521]), .C(poly13_shifted[507]), .D(n17755), .Z(n16241) );
  COND1XL U15708 ( .A(n17741), .B(n17491), .C(n16241), .Z(n10553) );
  CANR2XL U15709 ( .A(n17574), .B(Poly7[236]), .C(n17705), .D(
        poly7_shifted[236]), .Z(n16242) );
  COND1XL U15710 ( .A(n17087), .B(n17574), .C(n16242), .Z(n9868) );
  CANR2X1 U15711 ( .A(n17053), .B(Poly1[204]), .C(n18234), .D(
        poly1_shifted[204]), .Z(n16243) );
  COND1XL U15712 ( .A(n17087), .B(n17053), .C(n16243), .Z(n9153) );
  CANR2X1 U15713 ( .A(n12211), .B(poly2_shifted[24]), .C(n17523), .D(
        poly2_shifted[12]), .Z(n16244) );
  COND1XL U15714 ( .A(n17087), .B(n12211), .C(n16244), .Z(n8998) );
  CANR2X1 U15715 ( .A(n12977), .B(poly7_shifted[184]), .C(n17535), .D(
        poly7_shifted[172]), .Z(n16245) );
  COND1XL U15716 ( .A(n17087), .B(n12977), .C(n16245), .Z(n9932) );
  CANR2X1 U15717 ( .A(n12012), .B(poly1_shifted[87]), .C(n17998), .D(
        poly1_shifted[76]), .Z(n16246) );
  COND1XL U15718 ( .A(n17087), .B(n12012), .C(n16246), .Z(n9281) );
  CANR2X1 U15719 ( .A(n16425), .B(poly1_shifted[119]), .C(n17655), .D(
        poly1_shifted[108]), .Z(n16247) );
  COND1XL U15720 ( .A(n17087), .B(n16425), .C(n16247), .Z(n9249) );
  COND1XL U15721 ( .A(dataselector[61]), .B(n16249), .C(n16248), .Z(n16250) );
  CMXI2XL U15722 ( .A0(dataselector[15]), .A1(n16250), .S(n17831), .Z(n16251)
         );
  COND11XL U15723 ( .A(dataselector[8]), .B(n16252), .C(n17495), .D(n16251), 
        .Z(n8780) );
  CANR2XL U15724 ( .A(n18028), .B(poly7_shifted[306]), .C(n17215), .D(
        poly7_shifted[294]), .Z(n16253) );
  COND1XL U15725 ( .A(n17757), .B(n18028), .C(n16253), .Z(n9810) );
  CANR2X1 U15726 ( .A(n12009), .B(poly14_shifted[124]), .C(n17504), .D(
        poly14_shifted[108]), .Z(n16254) );
  COND1XL U15727 ( .A(n17087), .B(n12009), .C(n16254), .Z(n10297) );
  CANR2X1 U15728 ( .A(n12008), .B(poly14_shifted[156]), .C(n17508), .D(
        poly14_shifted[140]), .Z(n16255) );
  COND1XL U15729 ( .A(n17087), .B(n12008), .C(n16255), .Z(n10265) );
  CANR2X1 U15730 ( .A(n17444), .B(Poly14[300]), .C(n16919), .D(
        poly14_shifted[300]), .Z(n16256) );
  COND1XL U15731 ( .A(n17087), .B(n17444), .C(n16256), .Z(n10105) );
  CANR2X1 U15732 ( .A(n12175), .B(Poly8[12]), .C(n17620), .D(Poly8[94]), .Z(
        n16257) );
  COND1XL U15733 ( .A(n17087), .B(n12175), .C(n16257), .Z(n11389) );
  CENX1 U15734 ( .A(Poly2[68]), .B(Poly2[32]), .Z(n16258) );
  CENX1 U15735 ( .A(n17738), .B(n16258), .Z(n16259) );
  CNR2XL U15736 ( .A(n16259), .B(n17829), .Z(n16260) );
  CANR1XL U15737 ( .A(poly2_shifted[56]), .B(n17306), .C(n16260), .Z(n16261)
         );
  COND1XL U15738 ( .A(n17087), .B(n17306), .C(n16261), .Z(n8966) );
  CANR2X1 U15739 ( .A(n17525), .B(poly14_shifted[60]), .C(n17401), .D(
        poly14_shifted[44]), .Z(n16262) );
  COND1XL U15740 ( .A(n17087), .B(n17525), .C(n16262), .Z(n10361) );
  CANR2X1 U15741 ( .A(n18002), .B(poly14_shifted[28]), .C(n16702), .D(
        Poly14[297]), .Z(n16263) );
  COND1XL U15742 ( .A(n17087), .B(n18002), .C(n16263), .Z(n10393) );
  CANR2X1 U15743 ( .A(n13129), .B(Poly14[172]), .C(n17280), .D(
        poly14_shifted[172]), .Z(n16264) );
  COND1XL U15744 ( .A(n17087), .B(n13129), .C(n16264), .Z(n10233) );
  CANR2X1 U15745 ( .A(n12932), .B(poly14_shifted[284]), .C(n16919), .D(
        poly14_shifted[268]), .Z(n16265) );
  COND1XL U15746 ( .A(n17087), .B(n12932), .C(n16265), .Z(n10137) );
  CIVX2 U15747 ( .A(n18116), .Z(n16779) );
  CANR2X1 U15748 ( .A(n17525), .B(poly14_shifted[54]), .C(n17714), .D(
        poly14_shifted[38]), .Z(n16266) );
  COND1XL U15749 ( .A(n16779), .B(n17525), .C(n16266), .Z(n10367) );
  CANR2X1 U15750 ( .A(n13124), .B(poly13_shifted[20]), .C(n17504), .D(
        Poly13[520]), .Z(n16267) );
  COND1XL U15751 ( .A(n16779), .B(n13124), .C(n16267), .Z(n11054) );
  CANR2X1 U15752 ( .A(n13014), .B(Poly13[166]), .C(n16540), .D(
        poly13_shifted[166]), .Z(n16268) );
  COND1XL U15753 ( .A(n16779), .B(n13014), .C(n16268), .Z(n10894) );
  CANR2X1 U15754 ( .A(n17987), .B(poly13_shifted[436]), .C(n16702), .D(
        poly13_shifted[422]), .Z(n16269) );
  COND1XL U15755 ( .A(n16779), .B(n17987), .C(n16269), .Z(n10638) );
  CANR2X1 U15756 ( .A(n12008), .B(poly14_shifted[150]), .C(n17714), .D(
        poly14_shifted[134]), .Z(n16270) );
  COND1XL U15757 ( .A(n16779), .B(n12008), .C(n16270), .Z(n10271) );
  CANR2X1 U15758 ( .A(n13129), .B(Poly14[166]), .C(n17714), .D(
        poly14_shifted[166]), .Z(n16271) );
  COND1XL U15759 ( .A(n16779), .B(n13129), .C(n16271), .Z(n10239) );
  CNR2IXL U15760 ( .B(poly7_shifted[351]), .A(n17160), .Z(n16272) );
  CANR1XL U15761 ( .A(poly7_shifted[363]), .B(n13040), .C(n16272), .Z(n16273)
         );
  COND1XL U15762 ( .A(n17188), .B(n13040), .C(n16273), .Z(n9753) );
  CIVXL U15763 ( .A(Poly0[116]), .Z(n16277) );
  CANR2X1 U15764 ( .A(n18082), .B(n16274), .C(n17375), .D(poly0_shifted[116]), 
        .Z(n16275) );
  COND1XL U15765 ( .A(n16277), .B(n16276), .C(n16275), .Z(n9461) );
  CANR2X1 U15766 ( .A(n17615), .B(poly13_shifted[314]), .C(n17298), .D(
        poly13_shifted[300]), .Z(n16278) );
  COND1XL U15767 ( .A(n17087), .B(n17615), .C(n16278), .Z(n10760) );
  CANR2X1 U15768 ( .A(n17615), .B(poly13_shifted[326]), .C(n17099), .D(
        poly13_shifted[312]), .Z(n16279) );
  COND1XL U15769 ( .A(n17721), .B(n17615), .C(n16279), .Z(n10748) );
  CANR2X1 U15770 ( .A(n17615), .B(poly13_shifted[312]), .C(n17158), .D(
        poly13_shifted[298]), .Z(n16280) );
  COND1XL U15771 ( .A(n12014), .B(n17615), .C(n16280), .Z(n10762) );
  CANR2X1 U15772 ( .A(n17615), .B(poly13_shifted[322]), .C(n18234), .D(
        poly13_shifted[308]), .Z(n16281) );
  COND1XL U15773 ( .A(n17707), .B(n17615), .C(n16281), .Z(n10752) );
  CANR2X1 U15774 ( .A(n17615), .B(poly13_shifted[311]), .C(n18017), .D(
        poly13_shifted[297]), .Z(n16282) );
  COND1XL U15775 ( .A(n12002), .B(n17615), .C(n16282), .Z(n10763) );
  CANR2X1 U15776 ( .A(n17615), .B(poly13_shifted[331]), .C(poly13_shifted[317]), .D(n16947), .Z(n16283) );
  COND1XL U15777 ( .A(n17185), .B(n17615), .C(n16283), .Z(n10743) );
  CEOXL U15778 ( .A(Poly13[525]), .B(Poly13[280]), .Z(n16284) );
  CANR2X1 U15779 ( .A(n17615), .B(poly13_shifted[308]), .C(n17527), .D(n16284), 
        .Z(n16285) );
  COND1XL U15780 ( .A(n16779), .B(n17615), .C(n16285), .Z(n10766) );
  CANR2X1 U15781 ( .A(n17615), .B(poly13_shifted[313]), .C(n17285), .D(
        poly13_shifted[299]), .Z(n16286) );
  COND1XL U15782 ( .A(n16994), .B(n17615), .C(n16286), .Z(n10761) );
  CIVX2 U15783 ( .A(n18048), .Z(n17173) );
  CANR2XL U15784 ( .A(n17471), .B(poly7_shifted[93]), .C(n17206), .D(
        poly7_shifted[81]), .Z(n16287) );
  COND1XL U15785 ( .A(n17173), .B(n17471), .C(n16287), .Z(n10023) );
  CANR2XL U15786 ( .A(n18028), .B(poly7_shifted[317]), .C(n17136), .D(
        poly7_shifted[305]), .Z(n16288) );
  COND1XL U15787 ( .A(n17173), .B(n18028), .C(n16288), .Z(n9799) );
  CANR2X1 U15788 ( .A(n12977), .B(poly7_shifted[189]), .C(n16479), .D(
        poly7_shifted[177]), .Z(n16289) );
  COND1XL U15789 ( .A(n17173), .B(n12977), .C(n16289), .Z(n9927) );
  CANR2X1 U15790 ( .A(n13040), .B(poly7_shifted[360]), .C(n17535), .D(
        poly7_shifted[348]), .Z(n16290) );
  COND1XL U15791 ( .A(n11978), .B(n13040), .C(n16290), .Z(n9756) );
  CANR2X1 U15792 ( .A(n13040), .B(poly7_shifted[347]), .C(n17266), .D(
        poly7_shifted[335]), .Z(n16291) );
  COND1XL U15793 ( .A(n17196), .B(n13040), .C(n16291), .Z(n9769) );
  CANR2X1 U15794 ( .A(n13040), .B(poly7_shifted[349]), .C(n17545), .D(
        poly7_shifted[337]), .Z(n16292) );
  COND1XL U15795 ( .A(n17076), .B(n13040), .C(n16292), .Z(n9767) );
  CANR2X1 U15796 ( .A(n13040), .B(poly7_shifted[337]), .C(n17535), .D(
        poly7_shifted[325]), .Z(n16293) );
  COND1XL U15797 ( .A(n11991), .B(n13040), .C(n16293), .Z(n9779) );
  CANR2X1 U15798 ( .A(n13040), .B(poly7_shifted[359]), .C(n17545), .D(
        poly7_shifted[347]), .Z(n16294) );
  COND1XL U15799 ( .A(n17741), .B(n13040), .C(n16294), .Z(n9757) );
  CANR2X1 U15800 ( .A(n12287), .B(poly8_shifted[75]), .C(n17121), .D(
        poly8_shifted[61]), .Z(n16295) );
  COND1XL U15801 ( .A(n17185), .B(n12287), .C(n16295), .Z(n11340) );
  CANR2X1 U15802 ( .A(n12287), .B(poly8_shifted[49]), .C(n16372), .D(
        poly8_shifted[35]), .Z(n16296) );
  COND1XL U15803 ( .A(n13275), .B(n12287), .C(n16296), .Z(n11366) );
  CANR2X1 U15804 ( .A(n12287), .B(poly8_shifted[63]), .C(n17705), .D(
        poly8_shifted[49]), .Z(n16297) );
  COND1XL U15805 ( .A(n17173), .B(n12287), .C(n16297), .Z(n11352) );
  CANR2X1 U15806 ( .A(n12287), .B(poly8_shifted[54]), .C(n18234), .D(
        poly8_shifted[40]), .Z(n16298) );
  COND1XL U15807 ( .A(n17163), .B(n12287), .C(n16298), .Z(n11361) );
  CANR2X1 U15808 ( .A(n12287), .B(poly8_shifted[73]), .C(n17538), .D(
        poly8_shifted[59]), .Z(n16299) );
  COND1XL U15809 ( .A(n17741), .B(n12287), .C(n16299), .Z(n11342) );
  CANR2X1 U15810 ( .A(n12287), .B(poly8_shifted[67]), .C(n17280), .D(
        poly8_shifted[53]), .Z(n16300) );
  COND1XL U15811 ( .A(n17036), .B(n12287), .C(n16300), .Z(n11348) );
  CANR2X1 U15812 ( .A(n12287), .B(poly8_shifted[59]), .C(n17198), .D(
        poly8_shifted[45]), .Z(n16301) );
  COND1XL U15813 ( .A(n17065), .B(n12287), .C(n16301), .Z(n11356) );
  CANR2X1 U15814 ( .A(n18002), .B(poly14_shifted[18]), .C(n17523), .D(
        Poly14[287]), .Z(n16302) );
  COND1XL U15815 ( .A(n16303), .B(n18002), .C(n16302), .Z(n10403) );
  CANR2X1 U15816 ( .A(n18002), .B(poly14_shifted[38]), .C(n17714), .D(
        poly14_shifted[22]), .Z(n16304) );
  COND1XL U15817 ( .A(n17001), .B(n18002), .C(n16304), .Z(n10383) );
  CANR2X1 U15818 ( .A(n18002), .B(poly14_shifted[40]), .C(n16787), .D(
        poly14_shifted[24]), .Z(n16305) );
  COND1XL U15819 ( .A(n16179), .B(n18002), .C(n16305), .Z(n10381) );
  CANR2X1 U15820 ( .A(n18002), .B(poly14_shifted[30]), .C(n16307), .D(
        Poly14[299]), .Z(n16306) );
  COND1XL U15821 ( .A(n12764), .B(n18002), .C(n16306), .Z(n10391) );
  CANR2X1 U15822 ( .A(n18002), .B(poly14_shifted[46]), .C(n16307), .D(
        poly14_shifted[30]), .Z(n16308) );
  COND1XL U15823 ( .A(n13418), .B(n18002), .C(n16308), .Z(n10375) );
  CANR2X1 U15824 ( .A(n18002), .B(poly14_shifted[16]), .C(n18234), .D(
        Poly14[285]), .Z(n16309) );
  COND1XL U15825 ( .A(n12011), .B(n18002), .C(n16309), .Z(n10405) );
  CANR2XL U15826 ( .A(n18002), .B(poly14_shifted[32]), .C(n18017), .D(
        poly14_shifted[16]), .Z(n16310) );
  COND1XL U15827 ( .A(n17062), .B(n18002), .C(n16310), .Z(n10389) );
  CANR2X1 U15828 ( .A(n18002), .B(poly14_shifted[29]), .C(n17598), .D(
        Poly14[298]), .Z(n16311) );
  COND1XL U15829 ( .A(n17065), .B(n18002), .C(n16311), .Z(n10392) );
  CANR2X1 U15830 ( .A(n12192), .B(poly1_shifted[235]), .C(n16312), .D(
        poly1_shifted[224]), .Z(n16313) );
  COND1XL U15831 ( .A(n17751), .B(n12192), .C(n16313), .Z(n9133) );
  CANR2X1 U15832 ( .A(n12192), .B(poly1_shifted[259]), .C(n18047), .D(
        poly1_shifted[248]), .Z(n16314) );
  COND1XL U15833 ( .A(n17721), .B(n12192), .C(n16314), .Z(n9109) );
  CANR2XL U15834 ( .A(n17503), .B(Poly0[20]), .C(poly0_shifted[20]), .D(n18017), .Z(n16315) );
  COND1XL U15835 ( .A(n17506), .B(n16391), .C(n16315), .Z(n9557) );
  CANR2X1 U15836 ( .A(n12997), .B(poly12_shifted[19]), .C(n17655), .D(
        Poly12[114]), .Z(n16316) );
  COND1XL U15837 ( .A(n13275), .B(n12997), .C(n16316), .Z(n10529) );
  CANR2X1 U15838 ( .A(n12997), .B(poly12_shifted[17]), .C(n17655), .D(
        Poly12[112]), .Z(n16317) );
  COND1XL U15839 ( .A(n16950), .B(n12997), .C(n16317), .Z(n10531) );
  CANR2X1 U15840 ( .A(n16694), .B(poly14_shifted[257]), .C(n17655), .D(
        poly14_shifted[241]), .Z(n16318) );
  COND1XL U15841 ( .A(n17173), .B(n16694), .C(n16318), .Z(n10164) );
  CANR2X1 U15842 ( .A(n16694), .B(poly14_shifted[256]), .C(n17458), .D(
        poly14_shifted[240]), .Z(n16319) );
  COND1XL U15843 ( .A(n17211), .B(n16694), .C(n16319), .Z(n10165) );
  CANR2X1 U15844 ( .A(n16694), .B(poly14_shifted[271]), .C(n16323), .D(
        poly14_shifted[255]), .Z(n16320) );
  COND1XL U15845 ( .A(n17188), .B(n16694), .C(n16320), .Z(n10150) );
  CANR2X1 U15846 ( .A(n16694), .B(poly14_shifted[267]), .C(n17174), .D(
        poly14_shifted[251]), .Z(n16321) );
  COND1XL U15847 ( .A(n17741), .B(n16694), .C(n16321), .Z(n10154) );
  CANR2X1 U15848 ( .A(n16694), .B(poly14_shifted[264]), .C(n16427), .D(
        poly14_shifted[248]), .Z(n16322) );
  COND1XL U15849 ( .A(n17721), .B(n16694), .C(n16322), .Z(n10157) );
  CANR2X1 U15850 ( .A(n16694), .B(poly14_shifted[255]), .C(n16323), .D(
        poly14_shifted[239]), .Z(n16324) );
  COND1XL U15851 ( .A(n17196), .B(n16694), .C(n16324), .Z(n10166) );
  CANR2XL U15852 ( .A(n12900), .B(poly13_shifted[47]), .C(n17607), .D(
        poly13_shifted[33]), .Z(n16325) );
  COND1XL U15853 ( .A(n16950), .B(n12900), .C(n16325), .Z(n11027) );
  CANR2X1 U15854 ( .A(n18198), .B(poly1_shifted[302]), .C(n16326), .D(
        poly1_shifted[291]), .Z(n16327) );
  COND1XL U15855 ( .A(n13275), .B(n18198), .C(n16327), .Z(n9066) );
  CANR2X1 U15856 ( .A(n18198), .B(poly1_shifted[321]), .C(n17099), .D(
        poly1_shifted[310]), .Z(n16328) );
  COND1XL U15857 ( .A(n17753), .B(n18198), .C(n16328), .Z(n9047) );
  CANR2X1 U15858 ( .A(n18198), .B(poly1_shifted[323]), .C(n16644), .D(
        poly1_shifted[312]), .Z(n16329) );
  COND1XL U15859 ( .A(n17721), .B(n18198), .C(n16329), .Z(n9045) );
  CANR2X1 U15860 ( .A(n17471), .B(poly7_shifted[106]), .C(n17466), .D(
        poly7_shifted[94]), .Z(n16330) );
  COND1XL U15861 ( .A(n13418), .B(n17471), .C(n16330), .Z(n10010) );
  CANR2X1 U15862 ( .A(n17471), .B(poly7_shifted[107]), .C(n17290), .D(
        poly7_shifted[95]), .Z(n16331) );
  COND1XL U15863 ( .A(n17188), .B(n17471), .C(n16331), .Z(n10009) );
  CANR2X1 U15864 ( .A(n17471), .B(poly7_shifted[103]), .C(n17094), .D(
        poly7_shifted[91]), .Z(n16332) );
  COND1XL U15865 ( .A(n17741), .B(n17471), .C(n16332), .Z(n10013) );
  CANR2X1 U15866 ( .A(n17471), .B(poly7_shifted[85]), .C(n17198), .D(
        poly7_shifted[73]), .Z(n16333) );
  COND1XL U15867 ( .A(n17208), .B(n17471), .C(n16333), .Z(n10031) );
  CANR2X1 U15868 ( .A(n17471), .B(poly7_shifted[88]), .C(n17352), .D(
        poly7_shifted[76]), .Z(n16334) );
  COND1XL U15869 ( .A(n17087), .B(n17471), .C(n16334), .Z(n10028) );
  CANR2X1 U15870 ( .A(n12287), .B(poly8_shifted[56]), .C(n17535), .D(
        poly8_shifted[42]), .Z(n16335) );
  COND1XL U15871 ( .A(n12014), .B(n12287), .C(n16335), .Z(n11359) );
  CANR2X1 U15872 ( .A(n17471), .B(poly7_shifted[89]), .C(n17099), .D(
        poly7_shifted[77]), .Z(n16336) );
  COND1XL U15873 ( .A(n17090), .B(n17471), .C(n16336), .Z(n10027) );
  CANR2X1 U15874 ( .A(n12287), .B(poly8_shifted[68]), .C(n17755), .D(
        poly8_shifted[54]), .Z(n16337) );
  COND1XL U15875 ( .A(n17001), .B(n12287), .C(n16337), .Z(n11347) );
  CANR2X1 U15876 ( .A(n17471), .B(poly7_shifted[100]), .C(n17352), .D(
        poly7_shifted[88]), .Z(n16338) );
  COND1XL U15877 ( .A(n16179), .B(n17471), .C(n16338), .Z(n10016) );
  CANR2X1 U15878 ( .A(n17471), .B(poly7_shifted[87]), .C(n17458), .D(
        poly7_shifted[75]), .Z(n16339) );
  COND1XL U15879 ( .A(n16994), .B(n17471), .C(n16339), .Z(n10029) );
  CANR2X1 U15880 ( .A(n12287), .B(poly8_shifted[57]), .C(n17466), .D(
        poly8_shifted[43]), .Z(n16340) );
  COND1XL U15881 ( .A(n16605), .B(n12287), .C(n16340), .Z(n11358) );
  CANR2X1 U15882 ( .A(n12287), .B(poly8_shifted[62]), .C(n17705), .D(
        poly8_shifted[48]), .Z(n16341) );
  COND1XL U15883 ( .A(n17062), .B(n12287), .C(n16341), .Z(n11353) );
  CANR2X1 U15884 ( .A(n12287), .B(poly8_shifted[74]), .C(n17449), .D(
        poly8_shifted[60]), .Z(n16342) );
  COND1XL U15885 ( .A(n11978), .B(n12287), .C(n16342), .Z(n11341) );
  CANR2X1 U15886 ( .A(n17471), .B(poly7_shifted[90]), .C(n17533), .D(
        poly7_shifted[78]), .Z(n16343) );
  COND1XL U15887 ( .A(n12764), .B(n17471), .C(n16343), .Z(n10026) );
  CANR2X1 U15888 ( .A(n12287), .B(poly8_shifted[76]), .C(n17094), .D(
        poly8_shifted[62]), .Z(n16344) );
  COND1XL U15889 ( .A(n13418), .B(n12287), .C(n16344), .Z(n11339) );
  CANR2X1 U15890 ( .A(n17969), .B(poly13_shifted[80]), .C(n17390), .D(
        poly13_shifted[66]), .Z(n16345) );
  COND1XL U15891 ( .A(n16303), .B(n17969), .C(n16345), .Z(n10994) );
  CANR2X1 U15892 ( .A(n17969), .B(poly13_shifted[85]), .C(n17613), .D(
        poly13_shifted[71]), .Z(n16346) );
  COND1XL U15893 ( .A(n16939), .B(n17969), .C(n16346), .Z(n10989) );
  CANR2X1 U15894 ( .A(n17969), .B(poly13_shifted[83]), .C(n17705), .D(
        poly13_shifted[69]), .Z(n16347) );
  COND1XL U15895 ( .A(n11983), .B(n17969), .C(n16347), .Z(n10991) );
  CANR2X1 U15896 ( .A(n17491), .B(poly13_shifted[496]), .C(n17560), .D(
        poly13_shifted[482]), .Z(n16348) );
  COND1XL U15897 ( .A(n16303), .B(n17491), .C(n16348), .Z(n10578) );
  CIVX1 U15898 ( .A(dataselector[34]), .Z(n18237) );
  COND1XL U15899 ( .A(dataselector[34]), .B(n16349), .C(n12002), .Z(n16351) );
  CMXI2X1 U15900 ( .A0(n16351), .A1(dataselector[41]), .S(n16350), .Z(n16352)
         );
  COND11XL U15901 ( .A(dataselector[57]), .B(n17959), .C(n18237), .D(n16352), 
        .Z(n8754) );
  CANR2X1 U15902 ( .A(n12202), .B(Poly14[198]), .C(n17714), .D(
        poly14_shifted[198]), .Z(n16353) );
  COND1XL U15903 ( .A(n17757), .B(n12202), .C(n16353), .Z(n10207) );
  CANR2X1 U15904 ( .A(n12202), .B(Poly14[204]), .C(n17714), .D(
        poly14_shifted[204]), .Z(n16354) );
  COND1XL U15905 ( .A(n17218), .B(n12202), .C(n16354), .Z(n10201) );
  CEOXL U15906 ( .A(Poly14[288]), .B(Poly14[196]), .Z(n16355) );
  CANR2X1 U15907 ( .A(n12202), .B(Poly14[212]), .C(n17398), .D(n16355), .Z(
        n16356) );
  COND1XL U15908 ( .A(n16391), .B(n12202), .C(n16356), .Z(n10193) );
  CANR2X1 U15909 ( .A(n12202), .B(Poly14[208]), .C(n18234), .D(
        poly14_shifted[208]), .Z(n16357) );
  COND1XL U15910 ( .A(n17211), .B(n12202), .C(n16357), .Z(n10197) );
  CANR2X1 U15911 ( .A(n12202), .B(Poly14[207]), .C(n17449), .D(
        poly14_shifted[207]), .Z(n16358) );
  COND1XL U15912 ( .A(n17196), .B(n12202), .C(n16358), .Z(n10198) );
  CANR2X1 U15913 ( .A(n12202), .B(Poly14[201]), .C(n16695), .D(
        poly14_shifted[201]), .Z(n16359) );
  COND1XL U15914 ( .A(n17208), .B(n12202), .C(n16359), .Z(n10204) );
  CANR2X1 U15915 ( .A(n12202), .B(Poly14[197]), .C(n16787), .D(
        poly14_shifted[197]), .Z(n16360) );
  COND1XL U15916 ( .A(n11985), .B(n12202), .C(n16360), .Z(n10208) );
  CANR2X1 U15917 ( .A(n12202), .B(Poly14[203]), .C(n17755), .D(
        poly14_shifted[203]), .Z(n16361) );
  COND1XL U15918 ( .A(n16605), .B(n12202), .C(n16361), .Z(n10202) );
  CANR2X1 U15919 ( .A(n12202), .B(Poly14[202]), .C(n16427), .D(
        poly14_shifted[202]), .Z(n16362) );
  COND1XL U15920 ( .A(n12014), .B(n12202), .C(n16362), .Z(n10203) );
  CENX1 U15921 ( .A(Poly14[205]), .B(Poly14[291]), .Z(n16363) );
  CENX1 U15922 ( .A(Poly14[297]), .B(n16363), .Z(n16364) );
  CANR2X1 U15923 ( .A(n12202), .B(poly14_shifted[237]), .C(n17755), .D(n16364), 
        .Z(n16365) );
  COND1XL U15924 ( .A(n17185), .B(n12202), .C(n16365), .Z(n10184) );
  CENX1 U15925 ( .A(Poly14[289]), .B(Poly14[295]), .Z(n16366) );
  CENX1 U15926 ( .A(Poly14[203]), .B(n16366), .Z(n16367) );
  CANR2X1 U15927 ( .A(n12202), .B(poly14_shifted[235]), .C(n17174), .D(n16367), 
        .Z(n16368) );
  COND1XL U15928 ( .A(n17741), .B(n12202), .C(n16368), .Z(n10186) );
  CANR2X1 U15929 ( .A(n17610), .B(Poly1[152]), .C(n17545), .D(
        poly1_shifted[152]), .Z(n16369) );
  COND1XL U15930 ( .A(n17721), .B(n17610), .C(n16369), .Z(n9205) );
  CANR2X1 U15931 ( .A(n17610), .B(Poly1[153]), .C(n17613), .D(
        poly1_shifted[153]), .Z(n16370) );
  COND1XL U15932 ( .A(n17123), .B(n17610), .C(n16370), .Z(n9204) );
  CANR2X1 U15933 ( .A(n17610), .B(Poly1[155]), .C(n16372), .D(
        poly1_shifted[155]), .Z(n16371) );
  COND1XL U15934 ( .A(n17741), .B(n17610), .C(n16371), .Z(n9202) );
  CANR2X1 U15935 ( .A(n17610), .B(poly1_shifted[144]), .C(n16372), .D(
        poly1_shifted[133]), .Z(n16373) );
  COND1XL U15936 ( .A(n11995), .B(n17610), .C(n16373), .Z(n9224) );
  CANR2X1 U15937 ( .A(n17610), .B(poly1_shifted[152]), .C(n17613), .D(
        poly1_shifted[141]), .Z(n16374) );
  COND1XL U15938 ( .A(n17090), .B(n17610), .C(n16374), .Z(n9216) );
  CANR2X1 U15939 ( .A(n17238), .B(poly0_shifted[52]), .C(poly0_shifted[70]), 
        .D(n17500), .Z(n16375) );
  COND1XL U15940 ( .A(n17502), .B(n16391), .C(n16375), .Z(n9525) );
  CANR2X1 U15941 ( .A(n17667), .B(poly13_shifted[222]), .C(n17620), .D(
        poly13_shifted[208]), .Z(n16376) );
  COND1XL U15942 ( .A(n17062), .B(n17667), .C(n16376), .Z(n10852) );
  CANR2X1 U15943 ( .A(n17667), .B(poly13_shifted[234]), .C(n17755), .D(
        poly13_shifted[220]), .Z(n16377) );
  COND1XL U15944 ( .A(n11978), .B(n17667), .C(n16377), .Z(n10840) );
  CANR2X1 U15945 ( .A(n17667), .B(poly13_shifted[236]), .C(n17508), .D(
        poly13_shifted[222]), .Z(n16378) );
  COND1XL U15946 ( .A(n13418), .B(n17667), .C(n16378), .Z(n10838) );
  CANR2X1 U15947 ( .A(n17667), .B(poly13_shifted[233]), .C(n17755), .D(
        poly13_shifted[219]), .Z(n16379) );
  COND1XL U15948 ( .A(n17741), .B(n17667), .C(n16379), .Z(n10841) );
  CEOX1 U15949 ( .A(n16380), .B(dataselector[4]), .Z(n16383) );
  CANR2X1 U15950 ( .A(n16381), .B(n17832), .C(dataselector[11]), .D(n16410), 
        .Z(n16382) );
  COND1XL U15951 ( .A(n17829), .B(n16383), .C(n16382), .Z(n8784) );
  CENX1 U15952 ( .A(n16385), .B(n16384), .Z(n17820) );
  CEOXL U15953 ( .A(Poly7[406]), .B(n17820), .Z(n16386) );
  CENX1 U15954 ( .A(dataselector[63]), .B(n16386), .Z(n16389) );
  CANR2X1 U15955 ( .A(n13428), .B(n17832), .C(dataselector[2]), .D(n16410), 
        .Z(n16388) );
  COND1XL U15956 ( .A(n17826), .B(n16389), .C(n16388), .Z(n8793) );
  CANR2X1 U15957 ( .A(n12977), .B(Poly7[180]), .C(n17072), .D(
        poly7_shifted[180]), .Z(n16390) );
  COND1XL U15958 ( .A(n16391), .B(n12977), .C(n16390), .Z(n9924) );
  CANR2X1 U15959 ( .A(n17667), .B(poly13_shifted[220]), .C(n17755), .D(
        poly13_shifted[206]), .Z(n16392) );
  COND1XL U15960 ( .A(n12764), .B(n17667), .C(n16392), .Z(n10854) );
  CANR2X1 U15961 ( .A(n17667), .B(poly13_shifted[219]), .C(n17755), .D(
        poly13_shifted[205]), .Z(n16393) );
  COND1XL U15962 ( .A(n17090), .B(n17667), .C(n16393), .Z(n10855) );
  CANR2X1 U15963 ( .A(n17667), .B(poly13_shifted[217]), .C(n17094), .D(
        poly13_shifted[203]), .Z(n16394) );
  COND1XL U15964 ( .A(n16994), .B(n17667), .C(n16394), .Z(n10857) );
  CANR2X1 U15965 ( .A(n17667), .B(poly13_shifted[213]), .C(n18234), .D(
        poly13_shifted[199]), .Z(n16395) );
  COND1XL U15966 ( .A(n16939), .B(n17667), .C(n16395), .Z(n10861) );
  CANR2X1 U15967 ( .A(n17667), .B(poly13_shifted[228]), .C(n16702), .D(
        poly13_shifted[214]), .Z(n16396) );
  COND1XL U15968 ( .A(n17753), .B(n17667), .C(n16396), .Z(n10846) );
  CANR2X1 U15969 ( .A(n17667), .B(poly13_shifted[218]), .C(n17285), .D(
        poly13_shifted[204]), .Z(n16397) );
  COND1XL U15970 ( .A(n17087), .B(n17667), .C(n16397), .Z(n10856) );
  CANR2X1 U15971 ( .A(n17667), .B(poly13_shifted[216]), .C(n17285), .D(
        poly13_shifted[202]), .Z(n16398) );
  COND1XL U15972 ( .A(n12014), .B(n17667), .C(n16398), .Z(n10858) );
  CANR2X1 U15973 ( .A(n17667), .B(poly13_shifted[215]), .C(n17634), .D(
        poly13_shifted[201]), .Z(n16399) );
  COND1XL U15974 ( .A(n17208), .B(n17667), .C(n16399), .Z(n10859) );
  CANR2X1 U15975 ( .A(n17610), .B(Poly1[159]), .C(n18234), .D(
        poly1_shifted[159]), .Z(n16400) );
  COND1XL U15976 ( .A(n17188), .B(n17610), .C(n16400), .Z(n9198) );
  CANR2X1 U15977 ( .A(n17610), .B(poly1_shifted[140]), .C(n16372), .D(
        poly1_shifted[129]), .Z(n16401) );
  COND1XL U15978 ( .A(n17697), .B(n17610), .C(n16401), .Z(n9228) );
  CANR2X1 U15979 ( .A(n17610), .B(poly1_shifted[153]), .C(n17280), .D(
        poly1_shifted[142]), .Z(n16402) );
  COND1XL U15980 ( .A(n17699), .B(n17610), .C(n16402), .Z(n9215) );
  CANR2X1 U15981 ( .A(n17610), .B(poly1_shifted[146]), .C(n16919), .D(
        poly1_shifted[135]), .Z(n16403) );
  COND1XL U15982 ( .A(n16939), .B(n17610), .C(n16403), .Z(n9222) );
  CANR2X1 U15983 ( .A(n17610), .B(poly1_shifted[150]), .C(n17705), .D(
        poly1_shifted[139]), .Z(n16404) );
  COND1XL U15984 ( .A(n16994), .B(n17610), .C(n16404), .Z(n9218) );
  CANR2X1 U15985 ( .A(n17610), .B(poly1_shifted[161]), .C(n17755), .D(
        poly1_shifted[150]), .Z(n16405) );
  COND1XL U15986 ( .A(n17753), .B(n17610), .C(n16405), .Z(n9207) );
  CANR2X1 U15987 ( .A(n17610), .B(poly1_shifted[141]), .C(n16479), .D(
        poly1_shifted[130]), .Z(n16406) );
  COND1XL U15988 ( .A(n16303), .B(n17610), .C(n16406), .Z(n9227) );
  CENX1 U15989 ( .A(Poly7[407]), .B(n16407), .Z(n16408) );
  CENX1 U15990 ( .A(n16409), .B(n16408), .Z(n16412) );
  CANR2X1 U15991 ( .A(n18053), .B(n17832), .C(dataselector[3]), .D(n16410), 
        .Z(n16411) );
  COND1XL U15992 ( .A(n16412), .B(n17495), .C(n16411), .Z(n8792) );
  CANR2X1 U15993 ( .A(n12161), .B(Poly12[64]), .C(n17640), .D(
        poly12_shifted[64]), .Z(n16413) );
  COND1XL U15994 ( .A(n17751), .B(n12161), .C(n16413), .Z(n10468) );
  CANR2X1 U15995 ( .A(n17444), .B(Poly14[294]), .C(n16999), .D(
        poly14_shifted[294]), .Z(n16414) );
  COND1XL U15996 ( .A(n16779), .B(n17444), .C(n16414), .Z(n10111) );
  CANR1XL U15997 ( .A(poly11_shifted[21]), .B(n12185), .C(n16415), .Z(n16416)
         );
  COND1XL U15998 ( .A(n16779), .B(n12185), .C(n16416), .Z(n11183) );
  CANR2X1 U15999 ( .A(n17491), .B(poly13_shifted[515]), .C(n18234), .D(
        poly13_shifted[501]), .Z(n16417) );
  COND1XL U16000 ( .A(n12006), .B(n17491), .C(n16417), .Z(n10559) );
  CANR2X1 U16001 ( .A(n16694), .B(poly14_shifted[261]), .C(n16435), .D(
        poly14_shifted[245]), .Z(n16418) );
  COND1XL U16002 ( .A(n12006), .B(n16694), .C(n16418), .Z(n10160) );
  CEOXL U16003 ( .A(Poly12[126]), .B(Poly12[37]), .Z(n16419) );
  CANR2X1 U16004 ( .A(n12598), .B(Poly12[53]), .C(n17634), .D(n16419), .Z(
        n16420) );
  COND1XL U16005 ( .A(n12006), .B(n12598), .C(n16420), .Z(n10479) );
  CEOXL U16006 ( .A(Poly3[39]), .B(Poly3[72]), .Z(n16421) );
  CENX1 U16007 ( .A(Poly3[78]), .B(n16421), .Z(n16422) );
  CNR2XL U16008 ( .A(n17829), .B(n16422), .Z(n16423) );
  CANR1XL U16009 ( .A(Poly3[53]), .B(n17262), .C(n16423), .Z(n16424) );
  COND1XL U16010 ( .A(n12006), .B(n17587), .C(n16424), .Z(n8887) );
  CANR2XL U16011 ( .A(n16425), .B(poly1_shifted[128]), .C(n17998), .D(
        poly1_shifted[117]), .Z(n16426) );
  COND1XL U16012 ( .A(n12006), .B(n16425), .C(n16426), .Z(n9240) );
  CANR2X1 U16013 ( .A(n12009), .B(poly14_shifted[133]), .C(n16427), .D(
        poly14_shifted[117]), .Z(n16428) );
  COND1XL U16014 ( .A(n12006), .B(n12009), .C(n16428), .Z(n10288) );
  CANR2X1 U16015 ( .A(n12900), .B(poly13_shifted[67]), .C(n17508), .D(
        poly13_shifted[53]), .Z(n16429) );
  COND1XL U16016 ( .A(n12006), .B(n12900), .C(n16429), .Z(n11007) );
  CEOXL U16017 ( .A(Poly14[285]), .B(Poly14[165]), .Z(n16430) );
  CANR2X1 U16018 ( .A(n13129), .B(poly14_shifted[197]), .C(n18234), .D(n16430), 
        .Z(n16431) );
  COND1XL U16019 ( .A(n12006), .B(n13129), .C(n16431), .Z(n10224) );
  CANR2X1 U16020 ( .A(n18198), .B(poly1_shifted[320]), .C(n16540), .D(
        poly1_shifted[309]), .Z(n16432) );
  COND1XL U16021 ( .A(n12006), .B(n18198), .C(n16432), .Z(n9048) );
  CANR2X1 U16022 ( .A(n12997), .B(Poly12[21]), .C(n17401), .D(
        poly12_shifted[21]), .Z(n16433) );
  COND1XL U16023 ( .A(n12006), .B(n12997), .C(n16433), .Z(n10511) );
  CANR2XL U16024 ( .A(n17667), .B(poly13_shifted[227]), .C(n18234), .D(
        poly13_shifted[213]), .Z(n16434) );
  COND1XL U16025 ( .A(n12006), .B(n17667), .C(n16434), .Z(n10847) );
  CANR2X1 U16026 ( .A(n12932), .B(poly14_shifted[293]), .C(n16435), .D(
        poly14_shifted[277]), .Z(n16436) );
  COND1XL U16027 ( .A(n12006), .B(n12932), .C(n16436), .Z(n10128) );
  CEOXL U16028 ( .A(Poly14[289]), .B(Poly14[197]), .Z(n16437) );
  CANR2X1 U16029 ( .A(n12202), .B(Poly14[213]), .C(n17174), .D(n16437), .Z(
        n16438) );
  COND1XL U16030 ( .A(n12006), .B(n12202), .C(n16438), .Z(n10192) );
  CANR2X1 U16031 ( .A(n17615), .B(poly13_shifted[323]), .C(n16435), .D(
        poly13_shifted[309]), .Z(n16439) );
  COND1XL U16032 ( .A(n12006), .B(n17615), .C(n16439), .Z(n10751) );
  CANR2X1 U16033 ( .A(n12211), .B(Poly2[21]), .C(n17375), .D(poly2_shifted[21]), .Z(n16440) );
  COND1XL U16034 ( .A(n12006), .B(n12211), .C(n16440), .Z(n8989) );
  CANR2X1 U16035 ( .A(n13124), .B(poly13_shifted[35]), .C(n17072), .D(
        poly13_shifted[21]), .Z(n16441) );
  COND1XL U16036 ( .A(n12006), .B(n13124), .C(n16441), .Z(n11039) );
  CAN2XL U16037 ( .A(n18017), .B(poly12_shifted[85]), .Z(n16442) );
  CANR1XL U16038 ( .A(Poly12[85]), .B(n12161), .C(n16442), .Z(n16443) );
  COND1XL U16039 ( .A(n12006), .B(n12161), .C(n16443), .Z(n10447) );
  CANR2X1 U16040 ( .A(n15737), .B(poly3_shifted[35]), .C(n17508), .D(
        poly3_shifted[21]), .Z(n16444) );
  COND1XL U16041 ( .A(n12006), .B(n15737), .C(n16444), .Z(n8919) );
  CANR2X1 U16042 ( .A(n12012), .B(poly1_shifted[96]), .C(n17998), .D(
        poly1_shifted[85]), .Z(n16445) );
  COND1XL U16043 ( .A(n12006), .B(n12012), .C(n16445), .Z(n9272) );
  CANR2X1 U16044 ( .A(n17987), .B(poly13_shifted[451]), .C(poly13_shifted[437]), .D(n17755), .Z(n16446) );
  COND1XL U16045 ( .A(n12006), .B(n17987), .C(n16446), .Z(n10623) );
  CANR2X1 U16046 ( .A(n17592), .B(Poly13[277]), .C(n16700), .D(
        poly13_shifted[277]), .Z(n16447) );
  COND1XL U16047 ( .A(n12006), .B(n17592), .C(n16447), .Z(n10783) );
  CEOXL U16048 ( .A(Poly13[518]), .B(Poly13[391]), .Z(n16448) );
  CANR2X1 U16049 ( .A(n17043), .B(poly13_shifted[419]), .C(n18234), .D(n16448), 
        .Z(n16449) );
  COND1XL U16050 ( .A(n12006), .B(n17043), .C(n16449), .Z(n10655) );
  CANR2X1 U16051 ( .A(n17525), .B(poly14_shifted[69]), .C(n17620), .D(
        poly14_shifted[53]), .Z(n16450) );
  COND1XL U16052 ( .A(n12006), .B(n17525), .C(n16450), .Z(n10352) );
  CEOXL U16053 ( .A(Poly13[526]), .B(Poly13[167]), .Z(n16451) );
  CANR2X1 U16054 ( .A(n13014), .B(poly13_shifted[195]), .C(n17198), .D(n16451), 
        .Z(n16452) );
  COND1XL U16055 ( .A(n12006), .B(n13014), .C(n16452), .Z(n10879) );
  CANR2X1 U16056 ( .A(n12625), .B(poly7_shifted[285]), .C(n17535), .D(
        poly7_shifted[273]), .Z(n16453) );
  COND1XL U16057 ( .A(n17173), .B(n12625), .C(n16453), .Z(n9831) );
  CANR2X1 U16058 ( .A(n12625), .B(poly7_shifted[273]), .C(n17535), .D(
        poly7_shifted[261]), .Z(n16454) );
  COND1XL U16059 ( .A(n11981), .B(n12625), .C(n16454), .Z(n9843) );
  CANR2X1 U16060 ( .A(n12625), .B(poly7_shifted[271]), .C(n17290), .D(
        poly7_shifted[259]), .Z(n16455) );
  COND1XL U16061 ( .A(n13275), .B(n12625), .C(n16455), .Z(n9845) );
  CANR2X1 U16062 ( .A(n12625), .B(poly7_shifted[270]), .C(n17523), .D(
        poly7_shifted[258]), .Z(n16456) );
  COND1XL U16063 ( .A(n16303), .B(n12625), .C(n16456), .Z(n9846) );
  CANR2X1 U16064 ( .A(n12625), .B(poly7_shifted[295]), .C(n17598), .D(
        poly7_shifted[283]), .Z(n16457) );
  COND1XL U16065 ( .A(n17741), .B(n12625), .C(n16457), .Z(n9821) );
  CANR2X1 U16066 ( .A(n12625), .B(poly7_shifted[283]), .C(n17598), .D(
        poly7_shifted[271]), .Z(n16458) );
  COND1XL U16067 ( .A(n17196), .B(n12625), .C(n16458), .Z(n9833) );
  CANR2X1 U16068 ( .A(n12625), .B(poly7_shifted[296]), .C(n17383), .D(
        poly7_shifted[284]), .Z(n16459) );
  COND1XL U16069 ( .A(n11978), .B(n12625), .C(n16459), .Z(n9820) );
  CANR2X1 U16070 ( .A(n18198), .B(poly1_shifted[300]), .C(n17755), .D(
        poly1_shifted[289]), .Z(n16460) );
  COND1XL U16071 ( .A(n17697), .B(n18198), .C(n16460), .Z(n9068) );
  CANR2X1 U16072 ( .A(n16425), .B(poly1_shifted[108]), .C(n17527), .D(
        poly1_shifted[97]), .Z(n16461) );
  COND1XL U16073 ( .A(n17697), .B(n16425), .C(n16461), .Z(n9260) );
  CANR2X1 U16074 ( .A(n12977), .B(poly7_shifted[173]), .C(n17533), .D(
        poly7_shifted[161]), .Z(n16462) );
  COND1XL U16075 ( .A(n16950), .B(n12977), .C(n16462), .Z(n9943) );
  CANR2X1 U16076 ( .A(n17977), .B(poly13_shifted[167]), .C(n17094), .D(
        poly13_shifted[153]), .Z(n16463) );
  COND1XL U16077 ( .A(n17200), .B(n17977), .C(n16463), .Z(n10907) );
  CANR2X1 U16078 ( .A(n17977), .B(poly13_shifted[166]), .C(n17655), .D(
        poly13_shifted[152]), .Z(n16464) );
  COND1XL U16079 ( .A(n17721), .B(n17977), .C(n16464), .Z(n10908) );
  CANR2X1 U16080 ( .A(n17977), .B(Poly13[157]), .C(n17705), .D(
        poly13_shifted[157]), .Z(n16465) );
  COND1XL U16081 ( .A(n17185), .B(n17977), .C(n16465), .Z(n10903) );
  CANR2X1 U16082 ( .A(n17977), .B(Poly13[156]), .C(n17504), .D(
        poly13_shifted[156]), .Z(n16466) );
  COND1XL U16083 ( .A(n11978), .B(n17977), .C(n16466), .Z(n10904) );
  CANR2X1 U16084 ( .A(n17977), .B(poly13_shifted[142]), .C(n17613), .D(
        poly13_shifted[128]), .Z(n16467) );
  COND1XL U16085 ( .A(n12011), .B(n17977), .C(n16467), .Z(n10932) );
  CANR2X1 U16086 ( .A(n17977), .B(poly13_shifted[151]), .C(n17642), .D(
        poly13_shifted[137]), .Z(n16468) );
  COND1XL U16087 ( .A(n12002), .B(n17977), .C(n16468), .Z(n10923) );
  CANR2X1 U16088 ( .A(n17977), .B(poly13_shifted[163]), .C(n17755), .D(
        poly13_shifted[149]), .Z(n16469) );
  COND1XL U16089 ( .A(n12006), .B(n17977), .C(n16469), .Z(n10911) );
  CANR2X1 U16090 ( .A(n17977), .B(poly13_shifted[162]), .C(n17755), .D(
        poly13_shifted[148]), .Z(n16470) );
  COND1XL U16091 ( .A(n17707), .B(n17977), .C(n16470), .Z(n10912) );
  CANR2X1 U16092 ( .A(n17977), .B(poly13_shifted[150]), .C(n17280), .D(
        poly13_shifted[136]), .Z(n16471) );
  COND1XL U16093 ( .A(n17163), .B(n17977), .C(n16471), .Z(n10924) );
  CANR2X1 U16094 ( .A(n17977), .B(poly13_shifted[155]), .C(n18234), .D(
        poly13_shifted[141]), .Z(n16472) );
  COND1XL U16095 ( .A(n17065), .B(n17977), .C(n16472), .Z(n10919) );
  CANR2X1 U16096 ( .A(n17977), .B(poly13_shifted[152]), .C(n17705), .D(
        poly13_shifted[138]), .Z(n16473) );
  COND1XL U16097 ( .A(n12014), .B(n17977), .C(n16473), .Z(n10922) );
  CANR2X1 U16098 ( .A(n17977), .B(poly13_shifted[164]), .C(n16919), .D(
        poly13_shifted[150]), .Z(n16474) );
  COND1XL U16099 ( .A(n17001), .B(n17977), .C(n16474), .Z(n10910) );
  CANR2XL U16100 ( .A(n17977), .B(poly13_shifted[143]), .C(n18017), .D(
        poly13_shifted[129]), .Z(n16475) );
  COND1XL U16101 ( .A(n16950), .B(n17977), .C(n16475), .Z(n10931) );
  CANR2X1 U16102 ( .A(n13070), .B(poly7_shifted[153]), .C(n16479), .D(
        poly7_shifted[141]), .Z(n16476) );
  COND1XL U16103 ( .A(n17065), .B(n13070), .C(n16476), .Z(n9963) );
  CANR2X1 U16104 ( .A(n13070), .B(poly7_shifted[141]), .C(n16479), .D(
        poly7_shifted[129]), .Z(n16477) );
  COND1XL U16105 ( .A(n17697), .B(n13070), .C(n16477), .Z(n9975) );
  CANR2X1 U16106 ( .A(n13070), .B(poly7_shifted[169]), .C(n17178), .D(
        poly7_shifted[157]), .Z(n16478) );
  COND1XL U16107 ( .A(n17185), .B(n13070), .C(n16478), .Z(n9947) );
  CANR2X1 U16108 ( .A(n13070), .B(poly7_shifted[165]), .C(n16479), .D(
        poly7_shifted[153]), .Z(n16480) );
  COND1XL U16109 ( .A(n17123), .B(n13070), .C(n16480), .Z(n9951) );
  CANR2X1 U16110 ( .A(n13070), .B(poly7_shifted[167]), .C(n17535), .D(
        poly7_shifted[155]), .Z(n16481) );
  COND1XL U16111 ( .A(n17741), .B(n13070), .C(n16481), .Z(n9949) );
  CANR2X1 U16112 ( .A(n13070), .B(poly7_shifted[156]), .C(n17285), .D(
        poly7_shifted[144]), .Z(n16482) );
  COND1XL U16113 ( .A(n17211), .B(n13070), .C(n16482), .Z(n9960) );
  CEOXL U16114 ( .A(n17233), .B(Poly11[37]), .Z(n16483) );
  CANR2X1 U16115 ( .A(n17683), .B(Poly11[52]), .C(n18234), .D(n16483), .Z(
        n16484) );
  COND1XL U16116 ( .A(n17707), .B(n17747), .C(n16484), .Z(n11137) );
  CANR2X1 U16117 ( .A(n17525), .B(poly14_shifted[68]), .C(n17063), .D(
        poly14_shifted[52]), .Z(n16485) );
  COND1XL U16118 ( .A(n17707), .B(n17525), .C(n16485), .Z(n10353) );
  CANR2X1 U16119 ( .A(n17667), .B(poly13_shifted[226]), .C(n17705), .D(
        poly13_shifted[212]), .Z(n16486) );
  COND1XL U16120 ( .A(n17707), .B(n17667), .C(n16486), .Z(n10848) );
  CANR2X1 U16121 ( .A(n17955), .B(Poly9[84]), .C(n17466), .D(poly9_shifted[84]), .Z(n16487) );
  COND1XL U16122 ( .A(n17707), .B(n17955), .C(n16487), .Z(n11221) );
  CANR2X1 U16123 ( .A(n17574), .B(Poly7[244]), .C(n16488), .D(
        poly7_shifted[244]), .Z(n16489) );
  COND1XL U16124 ( .A(n17707), .B(n17574), .C(n16489), .Z(n9860) );
  CEOXL U16125 ( .A(Poly13[525]), .B(Poly13[166]), .Z(n16490) );
  CANR2X1 U16126 ( .A(n13014), .B(poly13_shifted[194]), .C(n17178), .D(n16490), 
        .Z(n16491) );
  COND1XL U16127 ( .A(n17707), .B(n13014), .C(n16491), .Z(n10880) );
  CANR2X1 U16128 ( .A(n17610), .B(poly1_shifted[159]), .C(n17280), .D(
        poly1_shifted[148]), .Z(n16492) );
  COND1XL U16129 ( .A(n17707), .B(n17610), .C(n16492), .Z(n9209) );
  CANR2X1 U16130 ( .A(n17491), .B(poly13_shifted[514]), .C(n17655), .D(
        poly13_shifted[500]), .Z(n16493) );
  COND1XL U16131 ( .A(n17707), .B(n17491), .C(n16493), .Z(n10560) );
  CANR2X1 U16132 ( .A(n16425), .B(poly1_shifted[127]), .C(n17343), .D(
        poly1_shifted[116]), .Z(n16494) );
  COND1XL U16133 ( .A(n17707), .B(n16425), .C(n16494), .Z(n9241) );
  CANR2XL U16134 ( .A(n12012), .B(poly1_shifted[95]), .C(poly1_shifted[84]), 
        .D(n18017), .Z(n16495) );
  COND1XL U16135 ( .A(n17707), .B(n12012), .C(n16495), .Z(n9273) );
  CANR2X1 U16136 ( .A(n17974), .B(poly13_shifted[130]), .C(n17755), .D(
        poly13_shifted[116]), .Z(n16496) );
  COND1XL U16137 ( .A(n17707), .B(n17974), .C(n16496), .Z(n10944) );
  CANR2X1 U16138 ( .A(n17731), .B(Poly9[20]), .C(n16695), .D(poly9_shifted[20]), .Z(n16497) );
  COND1XL U16139 ( .A(n17707), .B(n17731), .C(n16497), .Z(n11285) );
  CANR2X1 U16140 ( .A(n12210), .B(poly1_shifted[191]), .C(n17156), .D(
        poly1_shifted[180]), .Z(n16498) );
  COND1XL U16141 ( .A(n17707), .B(n12210), .C(n16498), .Z(n9177) );
  CANR2X1 U16142 ( .A(n12185), .B(Poly11[20]), .C(n18234), .D(
        poly11_shifted[20]), .Z(n16499) );
  COND1XL U16143 ( .A(n17707), .B(n12185), .C(n16499), .Z(n11169) );
  CANR2X1 U16144 ( .A(n18002), .B(poly14_shifted[36]), .C(n17613), .D(
        poly14_shifted[20]), .Z(n16500) );
  COND1XL U16145 ( .A(n16391), .B(n18002), .C(n16500), .Z(n10385) );
  CANR2X1 U16146 ( .A(n18191), .B(poly1_shifted[287]), .C(n17634), .D(
        poly1_shifted[276]), .Z(n16501) );
  COND1XL U16147 ( .A(n16391), .B(n18191), .C(n16501), .Z(n9081) );
  CANR2X1 U16148 ( .A(n18230), .B(Poly4[20]), .C(n16502), .D(poly4_shifted[20]), .Z(n16503) );
  COND1XL U16149 ( .A(n16391), .B(n18230), .C(n16503), .Z(n8836) );
  CANR2X1 U16150 ( .A(n12009), .B(poly14_shifted[132]), .C(n17504), .D(
        poly14_shifted[116]), .Z(n16504) );
  COND1XL U16151 ( .A(n16391), .B(n12009), .C(n16504), .Z(n10289) );
  CANR2X1 U16152 ( .A(n17273), .B(poly7_shifted[224]), .C(n17545), .D(
        poly7_shifted[212]), .Z(n16505) );
  COND1XL U16153 ( .A(n16391), .B(n17273), .C(n16505), .Z(n9892) );
  CANR2X1 U16154 ( .A(n13040), .B(poly7_shifted[352]), .C(n17072), .D(
        poly7_shifted[340]), .Z(n16506) );
  COND1XL U16155 ( .A(n16391), .B(n13040), .C(n16506), .Z(n9764) );
  CANR2XL U16156 ( .A(n12932), .B(poly14_shifted[292]), .C(n17206), .D(
        poly14_shifted[276]), .Z(n16507) );
  COND1XL U16157 ( .A(n16391), .B(n12932), .C(n16507), .Z(n10129) );
  CANR2X1 U16158 ( .A(n12211), .B(Poly2[20]), .C(n17203), .D(poly2_shifted[20]), .Z(n16508) );
  COND1XL U16159 ( .A(n16391), .B(n12211), .C(n16508), .Z(n8990) );
  CANR2XL U16160 ( .A(n18028), .B(poly7_shifted[320]), .C(n17206), .D(
        poly7_shifted[308]), .Z(n16509) );
  COND1XL U16161 ( .A(n16391), .B(n18028), .C(n16509), .Z(n9796) );
  CANR2X1 U16162 ( .A(n13070), .B(poly7_shifted[160]), .C(n17209), .D(
        poly7_shifted[148]), .Z(n16510) );
  COND1XL U16163 ( .A(n16391), .B(n13070), .C(n16510), .Z(n9956) );
  CANR2X1 U16164 ( .A(n12012), .B(poly1_shifted[103]), .C(n18234), .D(
        poly1_shifted[92]), .Z(n16511) );
  COND1XL U16165 ( .A(n11978), .B(n12012), .C(n16511), .Z(n9265) );
  CANR2X1 U16166 ( .A(n16425), .B(poly1_shifted[135]), .C(n17508), .D(
        poly1_shifted[124]), .Z(n16512) );
  COND1XL U16167 ( .A(n11978), .B(n16425), .C(n16512), .Z(n9233) );
  CANR2X1 U16168 ( .A(n17471), .B(poly7_shifted[104]), .C(n17449), .D(
        poly7_shifted[92]), .Z(n16513) );
  COND1XL U16169 ( .A(n11978), .B(n17471), .C(n16513), .Z(n10012) );
  CANR2X1 U16170 ( .A(n12977), .B(Poly7[188]), .C(n17401), .D(
        poly7_shifted[188]), .Z(n16514) );
  COND1XL U16171 ( .A(n11978), .B(n12977), .C(n16514), .Z(n9916) );
  CANR2XL U16172 ( .A(n18191), .B(poly1_shifted[295]), .C(n18234), .D(
        poly1_shifted[284]), .Z(n16515) );
  COND1XL U16173 ( .A(n11978), .B(n18191), .C(n16515), .Z(n9073) );
  CANR2X1 U16174 ( .A(n17266), .B(poly0_shifted[63]), .C(n17500), .D(
        poly0_shifted[81]), .Z(n16516) );
  COND1XL U16175 ( .A(n17502), .B(n17188), .C(n16516), .Z(n9514) );
  CANR2X1 U16176 ( .A(n17401), .B(poly0_shifted[55]), .C(n17500), .D(
        poly0_shifted[73]), .Z(n16517) );
  COND1XL U16177 ( .A(n17502), .B(n12296), .C(n16517), .Z(n9522) );
  CANR2X1 U16178 ( .A(n17613), .B(poly0_shifted[48]), .C(n17500), .D(
        poly0_shifted[66]), .Z(n16518) );
  COND1XL U16179 ( .A(n17502), .B(n17062), .C(n16518), .Z(n9529) );
  CANR2X1 U16180 ( .A(n17705), .B(poly0_shifted[60]), .C(n17500), .D(
        poly0_shifted[78]), .Z(n16519) );
  COND1XL U16181 ( .A(n17502), .B(n11978), .C(n16519), .Z(n9517) );
  CANR2X1 U16182 ( .A(n17266), .B(poly0_shifted[62]), .C(n17500), .D(
        poly0_shifted[80]), .Z(n16520) );
  COND1XL U16183 ( .A(n17502), .B(n17004), .C(n16520), .Z(n9515) );
  CANR2X1 U16184 ( .A(n17063), .B(poly0_shifted[47]), .C(n17500), .D(
        poly0_shifted[65]), .Z(n16521) );
  COND1XL U16185 ( .A(n17502), .B(n17196), .C(n16521), .Z(n9530) );
  CANR2X1 U16186 ( .A(n17655), .B(poly0_shifted[56]), .C(n17500), .D(
        poly0_shifted[74]), .Z(n16522) );
  COND1XL U16187 ( .A(n17502), .B(n17721), .C(n16522), .Z(n9521) );
  CANR2X1 U16188 ( .A(n17705), .B(poly0_shifted[53]), .C(n17500), .D(
        poly0_shifted[71]), .Z(n16523) );
  COND1XL U16189 ( .A(n17502), .B(n12006), .C(n16523), .Z(n9524) );
  CANR2X1 U16190 ( .A(n17655), .B(poly0_shifted[41]), .C(n17500), .D(
        poly0_shifted[59]), .Z(n16524) );
  COND1XL U16191 ( .A(n17502), .B(n17208), .C(n16524), .Z(n9536) );
  CANR2X1 U16192 ( .A(n18234), .B(poly0_shifted[42]), .C(n17500), .D(
        poly0_shifted[60]), .Z(n16525) );
  COND1XL U16193 ( .A(n17502), .B(n12014), .C(n16525), .Z(n9535) );
  CANR2X1 U16194 ( .A(n17613), .B(poly0_shifted[54]), .C(n17500), .D(
        poly0_shifted[72]), .Z(n16526) );
  COND1XL U16195 ( .A(n17502), .B(n17753), .C(n16526), .Z(n9523) );
  CANR2X1 U16196 ( .A(n17705), .B(poly0_shifted[61]), .C(n17500), .D(
        poly0_shifted[79]), .Z(n16527) );
  COND1XL U16197 ( .A(n17502), .B(n17185), .C(n16527), .Z(n9516) );
  CANR2X1 U16198 ( .A(n18047), .B(poly0_shifted[44]), .C(n17500), .D(
        poly0_shifted[62]), .Z(n16528) );
  COND1XL U16199 ( .A(n17502), .B(n17087), .C(n16528), .Z(n9533) );
  CANR2X1 U16200 ( .A(n17634), .B(poly0_shifted[49]), .C(n17500), .D(
        poly0_shifted[67]), .Z(n16529) );
  COND1XL U16201 ( .A(n17502), .B(n17076), .C(n16529), .Z(n9528) );
  CANR2X1 U16202 ( .A(n17203), .B(poly0_shifted[45]), .C(n17500), .D(
        poly0_shifted[63]), .Z(n16530) );
  COND1XL U16203 ( .A(n17502), .B(n17090), .C(n16530), .Z(n9532) );
  CANR2X1 U16204 ( .A(n17652), .B(Poly12[118]), .C(n17466), .D(
        poly12_shifted[118]), .Z(n16531) );
  COND1XL U16205 ( .A(n17753), .B(n17652), .C(n16531), .Z(n10414) );
  CANR2X1 U16206 ( .A(n17974), .B(poly13_shifted[118]), .C(n17508), .D(
        poly13_shifted[104]), .Z(n16532) );
  COND1XL U16207 ( .A(n17166), .B(n17974), .C(n16532), .Z(n10956) );
  CANR2X1 U16208 ( .A(n12900), .B(poly13_shifted[54]), .C(n17755), .D(
        poly13_shifted[40]), .Z(n16533) );
  COND1XL U16209 ( .A(n17166), .B(n12900), .C(n16533), .Z(n11020) );
  CANR2XL U16210 ( .A(n17471), .B(poly7_shifted[84]), .C(n17215), .D(
        poly7_shifted[72]), .Z(n16534) );
  COND1XL U16211 ( .A(n17166), .B(n17471), .C(n16534), .Z(n10032) );
  CANR2X1 U16212 ( .A(n13124), .B(poly13_shifted[22]), .C(n17634), .D(
        Poly13[522]), .Z(n16535) );
  COND1XL U16213 ( .A(n17166), .B(n13124), .C(n16535), .Z(n11052) );
  CANR2X1 U16214 ( .A(n12008), .B(poly14_shifted[152]), .C(n16540), .D(
        poly14_shifted[136]), .Z(n16536) );
  COND1XL U16215 ( .A(n17166), .B(n12008), .C(n16536), .Z(n10269) );
  CANR2X1 U16216 ( .A(n17982), .B(poly13_shifted[374]), .C(n17965), .D(
        poly13_shifted[360]), .Z(n16537) );
  COND1XL U16217 ( .A(n17166), .B(n17982), .C(n16537), .Z(n10700) );
  CANR2X1 U16218 ( .A(n17444), .B(Poly14[296]), .C(n16999), .D(
        poly14_shifted[296]), .Z(n16538) );
  COND1XL U16219 ( .A(n17166), .B(n17444), .C(n16538), .Z(n10109) );
  CANR2X1 U16220 ( .A(n13129), .B(Poly14[168]), .C(n16540), .D(
        poly14_shifted[168]), .Z(n16539) );
  COND1XL U16221 ( .A(n17166), .B(n13129), .C(n16539), .Z(n10237) );
  CANR2X1 U16222 ( .A(n12009), .B(poly14_shifted[120]), .C(n16540), .D(
        poly14_shifted[104]), .Z(n16541) );
  COND1XL U16223 ( .A(n17166), .B(n12009), .C(n16541), .Z(n10301) );
  CANR2X1 U16224 ( .A(n17430), .B(Poly13[520]), .C(n17504), .D(
        poly13_shifted[520]), .Z(n16542) );
  COND1XL U16225 ( .A(n17166), .B(n17430), .C(n16542), .Z(n10540) );
  CANR2X1 U16226 ( .A(n18018), .B(poly7_shifted[20]), .C(n17613), .D(
        Poly7[407]), .Z(n16543) );
  COND1XL U16227 ( .A(n17166), .B(n17564), .C(n16543), .Z(n10096) );
  CANR2X1 U16228 ( .A(n12977), .B(poly7_shifted[180]), .C(n17063), .D(
        poly7_shifted[168]), .Z(n16544) );
  COND1XL U16229 ( .A(n17166), .B(n12977), .C(n16544), .Z(n9936) );
  CANR2X1 U16230 ( .A(n17525), .B(poly14_shifted[56]), .C(n16787), .D(
        poly14_shifted[40]), .Z(n16545) );
  COND1XL U16231 ( .A(n17166), .B(n17525), .C(n16545), .Z(n10365) );
  CANR2X1 U16232 ( .A(n12625), .B(poly7_shifted[290]), .C(n17545), .D(
        poly7_shifted[278]), .Z(n16546) );
  COND1XL U16233 ( .A(n17001), .B(n12625), .C(n16546), .Z(n9826) );
  CANR2X1 U16234 ( .A(n12625), .B(poly7_shifted[289]), .C(n17613), .D(
        poly7_shifted[277]), .Z(n16547) );
  COND1XL U16235 ( .A(n12006), .B(n12625), .C(n16547), .Z(n9827) );
  CANR2X1 U16236 ( .A(n12625), .B(poly7_shifted[276]), .C(n17535), .D(
        poly7_shifted[264]), .Z(n16548) );
  COND1XL U16237 ( .A(n17166), .B(n12625), .C(n16548), .Z(n9840) );
  CANR2X1 U16238 ( .A(n12625), .B(poly7_shifted[288]), .C(n17535), .D(
        poly7_shifted[276]), .Z(n16549) );
  COND1XL U16239 ( .A(n16391), .B(n12625), .C(n16549), .Z(n9828) );
  CANR2X1 U16240 ( .A(n12625), .B(poly7_shifted[278]), .C(n17535), .D(
        poly7_shifted[266]), .Z(n16550) );
  COND1XL U16241 ( .A(n12014), .B(n12625), .C(n16550), .Z(n9838) );
  CANR2X1 U16242 ( .A(n12625), .B(poly7_shifted[280]), .C(n18047), .D(
        poly7_shifted[268]), .Z(n16551) );
  COND1XL U16243 ( .A(n17087), .B(n12625), .C(n16551), .Z(n9836) );
  CANR2X1 U16244 ( .A(n12625), .B(poly7_shifted[277]), .C(n17072), .D(
        poly7_shifted[265]), .Z(n16552) );
  COND1XL U16245 ( .A(n17208), .B(n12625), .C(n16552), .Z(n9839) );
  CANR2X1 U16246 ( .A(n12625), .B(poly7_shifted[299]), .C(n17642), .D(
        poly7_shifted[287]), .Z(n16553) );
  COND1XL U16247 ( .A(n17188), .B(n12625), .C(n16553), .Z(n9817) );
  CIVXL U16248 ( .A(poly15_shifted[57]), .Z(n16564) );
  CIVX1 U16249 ( .A(Poly15[53]), .Z(n16554) );
  CNR2X1 U16250 ( .A(Poly15[27]), .B(n16554), .Z(n16561) );
  CND2X1 U16251 ( .A(Poly15[27]), .B(n16554), .Z(n16559) );
  CNR2XL U16252 ( .A(n16555), .B(n16561), .Z(n16556) );
  CANR1XL U16253 ( .A(n16559), .B(n16556), .C(n12013), .Z(n16557) );
  CANR4CX1 U16254 ( .A(n16559), .B(n16558), .C(n16557), .D(n17376), .Z(n16560)
         );
  CANR2X1 U16255 ( .A(n17990), .B(poly13_shifted[486]), .C(n18047), .D(
        poly13_shifted[472]), .Z(n16566) );
  COND1XL U16256 ( .A(n17721), .B(n17990), .C(n16566), .Z(n10588) );
  CANR2X1 U16257 ( .A(n17595), .B(poly13_shifted[253]), .C(n17620), .D(
        poly13_shifted[239]), .Z(n16567) );
  COND1XL U16258 ( .A(n17196), .B(n17595), .C(n16567), .Z(n10821) );
  CANR2X1 U16259 ( .A(n17990), .B(poly13_shifted[472]), .C(n17755), .D(
        poly13_shifted[458]), .Z(n16568) );
  COND1XL U16260 ( .A(n12014), .B(n17990), .C(n16568), .Z(n10602) );
  CANR2XL U16261 ( .A(n17595), .B(poly13_shifted[239]), .C(poly13_shifted[225]), .D(n18017), .Z(n16569) );
  COND1XL U16262 ( .A(n16950), .B(n17595), .C(n16569), .Z(n10835) );
  CANR2X1 U16263 ( .A(n17595), .B(poly13_shifted[248]), .C(n17755), .D(
        poly13_shifted[234]), .Z(n16570) );
  COND1XL U16264 ( .A(n12014), .B(n17595), .C(n16570), .Z(n10826) );
  CANR2X1 U16265 ( .A(n17595), .B(poly13_shifted[250]), .C(n17705), .D(
        poly13_shifted[236]), .Z(n16571) );
  COND1XL U16266 ( .A(n17087), .B(n17595), .C(n16571), .Z(n10824) );
  CANR2X1 U16267 ( .A(n17595), .B(poly13_shifted[258]), .C(n17634), .D(
        poly13_shifted[244]), .Z(n16572) );
  COND1XL U16268 ( .A(n17707), .B(n17595), .C(n16572), .Z(n10816) );
  CANR2X1 U16269 ( .A(n17990), .B(poly13_shifted[487]), .C(n17613), .D(
        poly13_shifted[473]), .Z(n16573) );
  COND1XL U16270 ( .A(n17200), .B(n17990), .C(n16573), .Z(n10587) );
  CANR2X1 U16271 ( .A(n17595), .B(poly13_shifted[245]), .C(n17094), .D(
        poly13_shifted[231]), .Z(n16574) );
  COND1XL U16272 ( .A(n16939), .B(n17595), .C(n16574), .Z(n10829) );
  CANR2X1 U16273 ( .A(n17595), .B(poly13_shifted[268]), .C(n17538), .D(
        poly13_shifted[254]), .Z(n16575) );
  COND1XL U16274 ( .A(n13418), .B(n17595), .C(n16575), .Z(n10806) );
  CANR2X1 U16275 ( .A(n17595), .B(poly13_shifted[254]), .C(n17094), .D(
        poly13_shifted[240]), .Z(n16576) );
  COND1XL U16276 ( .A(n17062), .B(n17595), .C(n16576), .Z(n10820) );
  CANR2X1 U16277 ( .A(n17595), .B(poly13_shifted[240]), .C(n16702), .D(
        poly13_shifted[226]), .Z(n16577) );
  COND1XL U16278 ( .A(n16775), .B(n17595), .C(n16577), .Z(n10834) );
  CANR2X1 U16279 ( .A(n17595), .B(poly13_shifted[238]), .C(n17238), .D(
        poly13_shifted[224]), .Z(n16578) );
  COND1XL U16280 ( .A(n12011), .B(n17595), .C(n16578), .Z(n10836) );
  CANR2X1 U16281 ( .A(n17595), .B(poly13_shifted[263]), .C(n16700), .D(
        poly13_shifted[249]), .Z(n16579) );
  COND1XL U16282 ( .A(n17200), .B(n17595), .C(n16579), .Z(n10811) );
  CANR2X1 U16283 ( .A(n17595), .B(poly13_shifted[266]), .C(n17136), .D(
        poly13_shifted[252]), .Z(n16580) );
  COND1XL U16284 ( .A(n11978), .B(n17595), .C(n16580), .Z(n10808) );
  CANR2X1 U16285 ( .A(n17595), .B(poly13_shifted[241]), .C(n17466), .D(
        poly13_shifted[227]), .Z(n16581) );
  COND1XL U16286 ( .A(n13275), .B(n17595), .C(n16581), .Z(n10833) );
  CANR2XL U16287 ( .A(n17990), .B(poly13_shifted[462]), .C(n18017), .D(
        poly13_shifted[448]), .Z(n16582) );
  COND1XL U16288 ( .A(n12011), .B(n17990), .C(n16582), .Z(n10612) );
  CANR2X1 U16289 ( .A(n17990), .B(poly13_shifted[493]), .C(n16583), .D(
        poly13_shifted[479]), .Z(n16584) );
  COND1XL U16290 ( .A(n17188), .B(n17990), .C(n16584), .Z(n10581) );
  CANR2X1 U16291 ( .A(n17990), .B(poly13_shifted[482]), .C(n17072), .D(
        poly13_shifted[468]), .Z(n16585) );
  COND1XL U16292 ( .A(n17707), .B(n17990), .C(n16585), .Z(n10592) );
  CANR2X1 U16293 ( .A(n17990), .B(poly13_shifted[474]), .C(n17449), .D(
        poly13_shifted[460]), .Z(n16586) );
  COND1XL U16294 ( .A(n17218), .B(n17990), .C(n16586), .Z(n10600) );
  CANR2X1 U16295 ( .A(n17595), .B(poly13_shifted[246]), .C(n17285), .D(
        poly13_shifted[232]), .Z(n16587) );
  COND1XL U16296 ( .A(n17166), .B(n17595), .C(n16587), .Z(n10828) );
  CANR2X1 U16297 ( .A(n17990), .B(poly13_shifted[489]), .C(n17072), .D(
        poly13_shifted[475]), .Z(n16588) );
  COND1XL U16298 ( .A(n17741), .B(n17990), .C(n16588), .Z(n10585) );
  CANR2X1 U16299 ( .A(n17990), .B(poly13_shifted[490]), .C(n17356), .D(
        poly13_shifted[476]), .Z(n16589) );
  COND1XL U16300 ( .A(n11978), .B(n17990), .C(n16589), .Z(n10584) );
  CANR2X1 U16301 ( .A(n17595), .B(poly13_shifted[255]), .C(n17198), .D(
        poly13_shifted[241]), .Z(n16590) );
  COND1XL U16302 ( .A(n17076), .B(n17595), .C(n16590), .Z(n10819) );
  CANR2X1 U16303 ( .A(n17990), .B(poly13_shifted[475]), .C(n17998), .D(
        poly13_shifted[461]), .Z(n16591) );
  COND1XL U16304 ( .A(n17090), .B(n17990), .C(n16591), .Z(n10599) );
  CANR2X1 U16305 ( .A(n17990), .B(poly13_shifted[476]), .C(n16919), .D(
        poly13_shifted[462]), .Z(n16592) );
  COND1XL U16306 ( .A(n17699), .B(n17990), .C(n16592), .Z(n10598) );
  CANR2X1 U16307 ( .A(n12299), .B(poly1_shifted[57]), .C(n16435), .D(
        poly1_shifted[46]), .Z(n16593) );
  COND1XL U16308 ( .A(n17699), .B(n12299), .C(n16593), .Z(n9311) );
  CANR2X1 U16309 ( .A(n12299), .B(poly1_shifted[56]), .C(n17705), .D(
        poly1_shifted[45]), .Z(n16594) );
  COND1XL U16310 ( .A(n17090), .B(n12299), .C(n16594), .Z(n9312) );
  CANR2X1 U16311 ( .A(n12299), .B(Poly1[63]), .C(n18234), .D(poly1_shifted[63]), .Z(n16595) );
  COND1XL U16312 ( .A(n17188), .B(n12299), .C(n16595), .Z(n9294) );
  CANR2X1 U16313 ( .A(n12299), .B(Poly1[62]), .C(n17285), .D(poly1_shifted[62]), .Z(n16596) );
  COND1XL U16314 ( .A(n17004), .B(n12299), .C(n16596), .Z(n9295) );
  CANR2X1 U16315 ( .A(n12299), .B(Poly1[57]), .C(n18234), .D(poly1_shifted[57]), .Z(n16597) );
  COND1XL U16316 ( .A(n17123), .B(n12299), .C(n16597), .Z(n9300) );
  CANR2X1 U16317 ( .A(n12299), .B(Poly1[53]), .C(n17063), .D(poly1_shifted[53]), .Z(n16598) );
  COND1XL U16318 ( .A(n12006), .B(n12299), .C(n16598), .Z(n9304) );
  CANR2X1 U16319 ( .A(n12299), .B(Poly1[56]), .C(n17063), .D(poly1_shifted[56]), .Z(n16599) );
  COND1XL U16320 ( .A(n17721), .B(n12299), .C(n16599), .Z(n9301) );
  CANR2X1 U16321 ( .A(n12299), .B(Poly1[54]), .C(n17362), .D(poly1_shifted[54]), .Z(n16600) );
  COND1XL U16322 ( .A(n17753), .B(n12299), .C(n16600), .Z(n9303) );
  CANR2X1 U16323 ( .A(n12299), .B(poly1_shifted[63]), .C(n17401), .D(
        poly1_shifted[52]), .Z(n16601) );
  COND1XL U16324 ( .A(n16391), .B(n12299), .C(n16601), .Z(n9305) );
  CANR2X1 U16325 ( .A(n12299), .B(poly1_shifted[55]), .C(n17552), .D(
        poly1_shifted[44]), .Z(n16602) );
  COND1XL U16326 ( .A(n17087), .B(n12299), .C(n16602), .Z(n9313) );
  CANR2X1 U16327 ( .A(n17525), .B(poly14_shifted[75]), .C(n16999), .D(
        poly14_shifted[59]), .Z(n16603) );
  COND1XL U16328 ( .A(n17741), .B(n17525), .C(n16603), .Z(n10346) );
  CANR2X1 U16329 ( .A(n17525), .B(poly14_shifted[59]), .C(n16999), .D(
        poly14_shifted[43]), .Z(n16604) );
  COND1XL U16330 ( .A(n16605), .B(n17525), .C(n16604), .Z(n10362) );
  CANR2X1 U16331 ( .A(n17990), .B(poly13_shifted[492]), .C(n17504), .D(
        poly13_shifted[478]), .Z(n16606) );
  COND1XL U16332 ( .A(n13418), .B(n17990), .C(n16606), .Z(n10582) );
  CANR2X1 U16333 ( .A(n17990), .B(poly13_shifted[467]), .C(n17466), .D(
        poly13_shifted[453]), .Z(n16607) );
  COND1XL U16334 ( .A(n11985), .B(n17990), .C(n16607), .Z(n10607) );
  CANR2X1 U16335 ( .A(n17595), .B(poly13_shifted[260]), .C(n17285), .D(
        poly13_shifted[246]), .Z(n16608) );
  COND1XL U16336 ( .A(n17001), .B(n17595), .C(n16608), .Z(n10814) );
  CANR2X1 U16337 ( .A(n17990), .B(poly13_shifted[463]), .C(n17449), .D(
        poly13_shifted[449]), .Z(n16609) );
  COND1XL U16338 ( .A(n17697), .B(n17990), .C(n16609), .Z(n10611) );
  CANR2X1 U16339 ( .A(n17595), .B(poly13_shifted[259]), .C(n17094), .D(
        poly13_shifted[245]), .Z(n16610) );
  COND1XL U16340 ( .A(n12006), .B(n17595), .C(n16610), .Z(n10815) );
  CANR2X1 U16341 ( .A(n17969), .B(poly13_shifted[87]), .C(n17965), .D(
        poly13_shifted[73]), .Z(n16611) );
  COND1XL U16342 ( .A(n12002), .B(n17969), .C(n16611), .Z(n10987) );
  CANR2X1 U16343 ( .A(n17969), .B(poly13_shifted[108]), .C(n17280), .D(
        poly13_shifted[94]), .Z(n16612) );
  COND1XL U16344 ( .A(n13418), .B(n17969), .C(n16612), .Z(n10966) );
  CANR2X1 U16345 ( .A(n17969), .B(poly13_shifted[102]), .C(n17383), .D(
        poly13_shifted[88]), .Z(n16613) );
  COND1XL U16346 ( .A(n16179), .B(n17969), .C(n16613), .Z(n10972) );
  CANR2X1 U16347 ( .A(n17969), .B(poly13_shifted[94]), .C(n17280), .D(
        poly13_shifted[80]), .Z(n16614) );
  COND1XL U16348 ( .A(n17062), .B(n17969), .C(n16614), .Z(n10980) );
  CANR2X1 U16349 ( .A(n17969), .B(poly13_shifted[78]), .C(n17634), .D(
        poly13_shifted[64]), .Z(n16615) );
  COND1XL U16350 ( .A(n17751), .B(n17969), .C(n16615), .Z(n10996) );
  CANR2X1 U16351 ( .A(n17969), .B(poly13_shifted[106]), .C(n17755), .D(
        poly13_shifted[92]), .Z(n16616) );
  COND1XL U16352 ( .A(n11978), .B(n17969), .C(n16616), .Z(n10968) );
  CANR2XL U16353 ( .A(n17969), .B(poly13_shifted[99]), .C(n18017), .D(
        poly13_shifted[85]), .Z(n16617) );
  COND1XL U16354 ( .A(n12006), .B(n17969), .C(n16617), .Z(n10975) );
  CANR2X1 U16355 ( .A(n13070), .B(poly7_shifted[168]), .C(n17998), .D(
        poly7_shifted[156]), .Z(n16618) );
  COND1XL U16356 ( .A(n11978), .B(n13070), .C(n16618), .Z(n9948) );
  CANR2X1 U16357 ( .A(n13070), .B(poly7_shifted[151]), .C(n18234), .D(
        poly7_shifted[139]), .Z(n16619) );
  COND1XL U16358 ( .A(n16994), .B(n13070), .C(n16619), .Z(n9965) );
  CANR2X1 U16359 ( .A(n13070), .B(poly7_shifted[152]), .C(n17362), .D(
        poly7_shifted[140]), .Z(n16620) );
  COND1XL U16360 ( .A(n17087), .B(n13070), .C(n16620), .Z(n9964) );
  CANR2X1 U16361 ( .A(n13070), .B(poly7_shifted[161]), .C(n17533), .D(
        poly7_shifted[149]), .Z(n16621) );
  COND1XL U16362 ( .A(n12006), .B(n13070), .C(n16621), .Z(n9955) );
  CANR2X1 U16363 ( .A(n13070), .B(poly7_shifted[154]), .C(n16427), .D(
        poly7_shifted[142]), .Z(n16622) );
  COND1XL U16364 ( .A(n12764), .B(n13070), .C(n16622), .Z(n9962) );
  CANR2X1 U16365 ( .A(n13070), .B(poly7_shifted[140]), .C(n17466), .D(
        poly7_shifted[128]), .Z(n16623) );
  COND1XL U16366 ( .A(n12011), .B(n13070), .C(n16623), .Z(n9976) );
  CANR2X1 U16367 ( .A(n13070), .B(poly7_shifted[162]), .C(n16695), .D(
        poly7_shifted[150]), .Z(n16624) );
  COND1XL U16368 ( .A(n17753), .B(n13070), .C(n16624), .Z(n9954) );
  CANR2X1 U16369 ( .A(n13070), .B(poly7_shifted[164]), .C(n17552), .D(
        poly7_shifted[152]), .Z(n16625) );
  COND1XL U16370 ( .A(n17721), .B(n13070), .C(n16625), .Z(n9952) );
  CANR2X1 U16371 ( .A(n13070), .B(poly7_shifted[142]), .C(n17266), .D(
        poly7_shifted[130]), .Z(n16626) );
  COND1XL U16372 ( .A(n16775), .B(n13070), .C(n16626), .Z(n9974) );
  CANR2X1 U16373 ( .A(n13070), .B(poly7_shifted[149]), .C(n17094), .D(
        poly7_shifted[137]), .Z(n16627) );
  COND1XL U16374 ( .A(n17208), .B(n13070), .C(n16627), .Z(n9967) );
  CANR2X1 U16375 ( .A(n17592), .B(Poly13[281]), .C(n17072), .D(
        poly13_shifted[281]), .Z(n16628) );
  COND1XL U16376 ( .A(n17200), .B(n17592), .C(n16628), .Z(n10779) );
  CEOXL U16377 ( .A(Poly13[514]), .B(Poly13[269]), .Z(n16629) );
  CANR2X1 U16378 ( .A(n17592), .B(poly13_shifted[297]), .C(n17458), .D(n16629), 
        .Z(n16630) );
  COND1XL U16379 ( .A(n17741), .B(n17592), .C(n16630), .Z(n10777) );
  CANR2XL U16380 ( .A(n17592), .B(poly13_shifted[278]), .C(poly13_shifted[264]), .D(n18017), .Z(n16631) );
  COND1XL U16381 ( .A(n17163), .B(n17592), .C(n16631), .Z(n10796) );
  CANR2X1 U16382 ( .A(n17592), .B(Poly13[278]), .C(n17705), .D(
        poly13_shifted[278]), .Z(n16632) );
  COND1XL U16383 ( .A(n17001), .B(n17592), .C(n16632), .Z(n10782) );
  CANR2X1 U16384 ( .A(n17652), .B(Poly12[96]), .C(n17655), .D(
        poly12_shifted[96]), .Z(n16633) );
  COND1XL U16385 ( .A(n17751), .B(n17652), .C(n16633), .Z(n10436) );
  CANR2X1 U16386 ( .A(n17652), .B(Poly12[116]), .C(n17401), .D(
        poly12_shifted[116]), .Z(n16634) );
  COND1XL U16387 ( .A(n17707), .B(n17652), .C(n16634), .Z(n10416) );
  CANR2X1 U16388 ( .A(n17652), .B(Poly12[117]), .C(n17613), .D(
        poly12_shifted[117]), .Z(n16635) );
  COND1XL U16389 ( .A(n12006), .B(n17652), .C(n16635), .Z(n10415) );
  CANR2X1 U16390 ( .A(n17652), .B(Poly12[121]), .C(n16479), .D(
        poly12_shifted[121]), .Z(n16636) );
  COND1XL U16391 ( .A(n17123), .B(n17652), .C(n16636), .Z(n10411) );
  CANR2X1 U16392 ( .A(n17652), .B(Poly12[120]), .C(n17613), .D(
        poly12_shifted[120]), .Z(n16637) );
  COND1XL U16393 ( .A(n17721), .B(n17652), .C(n16637), .Z(n10412) );
  CANR2X1 U16394 ( .A(n17652), .B(Poly12[113]), .C(n17356), .D(
        poly12_shifted[113]), .Z(n16638) );
  COND1XL U16395 ( .A(n17173), .B(n17652), .C(n16638), .Z(n10419) );
  CANR2X1 U16396 ( .A(n17652), .B(Poly12[125]), .C(n17508), .D(
        poly12_shifted[125]), .Z(n16639) );
  COND1XL U16397 ( .A(n17185), .B(n17652), .C(n16639), .Z(n10407) );
  CANR2XL U16398 ( .A(n17652), .B(Poly12[123]), .C(n18017), .D(
        poly12_shifted[123]), .Z(n16640) );
  COND1XL U16399 ( .A(n17741), .B(n17652), .C(n16640), .Z(n10409) );
  CANR2X1 U16400 ( .A(n12625), .B(poly7_shifted[298]), .C(n16307), .D(
        poly7_shifted[286]), .Z(n16641) );
  COND1XL U16401 ( .A(n13418), .B(n12625), .C(n16641), .Z(n9818) );
  CANR2X1 U16402 ( .A(n12625), .B(poly7_shifted[274]), .C(n16583), .D(
        poly7_shifted[262]), .Z(n16642) );
  COND1XL U16403 ( .A(n17757), .B(n12625), .C(n16642), .Z(n9842) );
  CANR2X1 U16404 ( .A(n12625), .B(poly7_shifted[269]), .C(n16985), .D(
        poly7_shifted[257]), .Z(n16643) );
  COND1XL U16405 ( .A(n17697), .B(n12625), .C(n16643), .Z(n9847) );
  CANR2X1 U16406 ( .A(n12958), .B(poly14_shifted[110]), .C(n16644), .D(
        poly14_shifted[94]), .Z(n16645) );
  COND1XL U16407 ( .A(n13418), .B(n12958), .C(n16645), .Z(n10311) );
  CANR2X1 U16408 ( .A(n12958), .B(poly14_shifted[82]), .C(n17527), .D(
        poly14_shifted[66]), .Z(n16646) );
  COND1XL U16409 ( .A(n16775), .B(n12958), .C(n16646), .Z(n10339) );
  CANR2X1 U16410 ( .A(n12958), .B(poly14_shifted[104]), .C(n16787), .D(
        poly14_shifted[88]), .Z(n16647) );
  COND1XL U16411 ( .A(n16179), .B(n12958), .C(n16647), .Z(n10317) );
  CANR2X1 U16412 ( .A(n12262), .B(Poly9[112]), .C(n17755), .D(
        poly9_shifted[112]), .Z(n16648) );
  COND1XL U16413 ( .A(n17211), .B(n12262), .C(n16648), .Z(n11193) );
  CANR2X1 U16414 ( .A(n18018), .B(poly7_shifted[28]), .C(n17121), .D(
        poly7_shifted[16]), .Z(n16649) );
  COND1XL U16415 ( .A(n17211), .B(n18018), .C(n16649), .Z(n10088) );
  CANR2X1 U16416 ( .A(n12210), .B(poly1_shifted[187]), .C(n17121), .D(
        poly1_shifted[176]), .Z(n16650) );
  COND1XL U16417 ( .A(n17211), .B(n12210), .C(n16650), .Z(n9181) );
  CANR2X1 U16418 ( .A(n12625), .B(poly7_shifted[284]), .C(n17383), .D(
        poly7_shifted[272]), .Z(n16651) );
  COND1XL U16419 ( .A(n17211), .B(n12625), .C(n16651), .Z(n9832) );
  CANR2X1 U16420 ( .A(n12977), .B(poly7_shifted[188]), .C(n17642), .D(
        poly7_shifted[176]), .Z(n16652) );
  COND1XL U16421 ( .A(n17211), .B(n12977), .C(n16652), .Z(n9928) );
  CANR2X1 U16422 ( .A(n15737), .B(poly3_shifted[30]), .C(n17356), .D(
        poly3_shifted[16]), .Z(n16653) );
  COND1XL U16423 ( .A(n17211), .B(n15737), .C(n16653), .Z(n8924) );
  CANR2X1 U16424 ( .A(n17273), .B(poly7_shifted[220]), .C(n17288), .D(
        poly7_shifted[208]), .Z(n16654) );
  COND1XL U16425 ( .A(n17211), .B(n17273), .C(n16654), .Z(n9896) );
  CANR2X1 U16426 ( .A(n12185), .B(poly11_shifted[31]), .C(n17705), .D(
        poly11_shifted[16]), .Z(n16655) );
  COND1XL U16427 ( .A(n17211), .B(n12185), .C(n16655), .Z(n11173) );
  CANR2X1 U16428 ( .A(n12012), .B(poly1_shifted[91]), .C(n18234), .D(
        poly1_shifted[80]), .Z(n16656) );
  COND1XL U16429 ( .A(n17211), .B(n12012), .C(n16656), .Z(n9277) );
  CANR2X1 U16430 ( .A(n17471), .B(poly7_shifted[92]), .C(n17458), .D(
        poly7_shifted[80]), .Z(n16657) );
  COND1XL U16431 ( .A(n17211), .B(n17471), .C(n16657), .Z(n10024) );
  CANR2X1 U16432 ( .A(n17671), .B(poly0_shifted[159]), .C(n17063), .D(
        poly0_shifted[141]), .Z(n16658) );
  COND1XL U16433 ( .A(n17674), .B(n17090), .C(n16658), .Z(n9436) );
  CANR2X1 U16434 ( .A(n17671), .B(Poly0[152]), .C(n17375), .D(
        poly0_shifted[152]), .Z(n16659) );
  COND1XL U16435 ( .A(n17674), .B(n17721), .C(n16659), .Z(n9425) );
  CANR2X1 U16436 ( .A(n12900), .B(poly13_shifted[63]), .C(n17072), .D(
        poly13_shifted[49]), .Z(n16660) );
  COND1XL U16437 ( .A(n17173), .B(n12900), .C(n16660), .Z(n11011) );
  CANR2X1 U16438 ( .A(n17592), .B(Poly13[273]), .C(n17298), .D(
        poly13_shifted[273]), .Z(n16661) );
  COND1XL U16439 ( .A(n17173), .B(n17592), .C(n16661), .Z(n10787) );
  CANR2X1 U16440 ( .A(n17615), .B(poly13_shifted[319]), .C(n17755), .D(
        poly13_shifted[305]), .Z(n16662) );
  COND1XL U16441 ( .A(n17173), .B(n17615), .C(n16662), .Z(n10755) );
  CANR2X1 U16442 ( .A(n17969), .B(poly13_shifted[95]), .C(n18234), .D(
        poly13_shifted[81]), .Z(n16663) );
  COND1XL U16443 ( .A(n17173), .B(n17969), .C(n16663), .Z(n10979) );
  CANR2XL U16444 ( .A(n17332), .B(poly1_shifted[339]), .C(n18017), .D(
        poly1_shifted[328]), .Z(n16664) );
  COND1XL U16445 ( .A(n17163), .B(n17332), .C(n16664), .Z(n9029) );
  CANR2X1 U16446 ( .A(n17332), .B(poly1_shifted[337]), .C(n17545), .D(
        poly1_shifted[326]), .Z(n16665) );
  COND1XL U16447 ( .A(n17757), .B(n17332), .C(n16665), .Z(n9031) );
  CANR2X1 U16448 ( .A(n17332), .B(poly1_shifted[333]), .C(n18234), .D(
        poly1_shifted[322]), .Z(n16666) );
  COND1XL U16449 ( .A(n16303), .B(n17332), .C(n16666), .Z(n9035) );
  CANR2X1 U16450 ( .A(n17332), .B(poly1_shifted[334]), .C(n17209), .D(
        poly1_shifted[323]), .Z(n16667) );
  COND1XL U16451 ( .A(n13275), .B(n17332), .C(n16667), .Z(n9034) );
  CANR2X1 U16452 ( .A(n17332), .B(poly1_shifted[344]), .C(n17634), .D(
        poly1_shifted[333]), .Z(n16668) );
  COND1XL U16453 ( .A(n17090), .B(n17332), .C(n16668), .Z(n9024) );
  CANR2X1 U16454 ( .A(n17332), .B(poly1_shifted[332]), .C(n17552), .D(
        poly1_shifted[321]), .Z(n16669) );
  COND1XL U16455 ( .A(n17697), .B(n17332), .C(n16669), .Z(n9036) );
  CANR2X1 U16456 ( .A(n17332), .B(poly1_shifted[331]), .C(n17072), .D(
        poly1_shifted[320]), .Z(n16670) );
  COND1XL U16457 ( .A(n12011), .B(n17332), .C(n16670), .Z(n9037) );
  CANR2X1 U16458 ( .A(n17332), .B(Poly1[341]), .C(n17560), .D(
        poly1_shifted[341]), .Z(n16671) );
  COND1XL U16459 ( .A(n12006), .B(n17332), .C(n16671), .Z(n9016) );
  CANR2X1 U16460 ( .A(n17332), .B(poly1_shifted[346]), .C(n17642), .D(
        poly1_shifted[335]), .Z(n16672) );
  COND1XL U16461 ( .A(n17196), .B(n17332), .C(n16672), .Z(n9022) );
  CANR2X1 U16462 ( .A(n17987), .B(poly13_shifted[447]), .C(n17504), .D(
        poly13_shifted[433]), .Z(n16673) );
  COND1XL U16463 ( .A(n17173), .B(n17987), .C(n16673), .Z(n10627) );
  CANR2X1 U16464 ( .A(n17667), .B(poly13_shifted[223]), .C(n17640), .D(
        poly13_shifted[209]), .Z(n16674) );
  COND1XL U16465 ( .A(n17173), .B(n17667), .C(n16674), .Z(n10851) );
  CANR2X1 U16466 ( .A(n17977), .B(poly13_shifted[154]), .C(n17348), .D(
        poly13_shifted[140]), .Z(n16675) );
  COND1XL U16467 ( .A(n17218), .B(n17977), .C(n16675), .Z(n10920) );
  CANR2X1 U16468 ( .A(n17969), .B(poly13_shifted[91]), .C(n17642), .D(
        poly13_shifted[77]), .Z(n16676) );
  COND1XL U16469 ( .A(n17090), .B(n17969), .C(n16676), .Z(n10983) );
  CANR2X1 U16470 ( .A(n17969), .B(poly13_shifted[92]), .C(n17755), .D(
        poly13_shifted[78]), .Z(n16677) );
  COND1XL U16471 ( .A(n12764), .B(n17969), .C(n16677), .Z(n10982) );
  CANR2X1 U16472 ( .A(n17969), .B(poly13_shifted[103]), .C(n17156), .D(
        poly13_shifted[89]), .Z(n16678) );
  COND1XL U16473 ( .A(n17123), .B(n17969), .C(n16678), .Z(n10971) );
  CANR2XL U16474 ( .A(n17969), .B(poly13_shifted[88]), .C(poly13_shifted[74]), 
        .D(n18017), .Z(n16679) );
  COND1XL U16475 ( .A(n12014), .B(n17969), .C(n16679), .Z(n10986) );
  CANR2X1 U16476 ( .A(n17969), .B(poly13_shifted[105]), .C(n17642), .D(
        poly13_shifted[91]), .Z(n16680) );
  COND1XL U16477 ( .A(n17741), .B(n17969), .C(n16680), .Z(n10969) );
  CANR2X1 U16478 ( .A(n17969), .B(poly13_shifted[89]), .C(n17343), .D(
        poly13_shifted[75]), .Z(n16681) );
  COND1XL U16479 ( .A(n16994), .B(n17969), .C(n16681), .Z(n10985) );
  CANR2X1 U16480 ( .A(n17969), .B(poly13_shifted[98]), .C(n16323), .D(
        poly13_shifted[84]), .Z(n16682) );
  COND1XL U16481 ( .A(n16391), .B(n17969), .C(n16682), .Z(n10976) );
  CANR2X1 U16482 ( .A(n17969), .B(poly13_shifted[84]), .C(n16702), .D(
        poly13_shifted[70]), .Z(n16683) );
  COND1XL U16483 ( .A(n16779), .B(n17969), .C(n16683), .Z(n10990) );
  CANR2X1 U16484 ( .A(n17969), .B(poly13_shifted[90]), .C(n17266), .D(
        poly13_shifted[76]), .Z(n16684) );
  COND1XL U16485 ( .A(n17087), .B(n17969), .C(n16684), .Z(n10984) );
  CANR2X1 U16486 ( .A(n16694), .B(poly14_shifted[269]), .C(n17755), .D(
        poly14_shifted[253]), .Z(n16685) );
  COND1XL U16487 ( .A(n17185), .B(n16694), .C(n16685), .Z(n10152) );
  CANR2X1 U16488 ( .A(n16694), .B(poly14_shifted[268]), .C(n16919), .D(
        poly14_shifted[252]), .Z(n16686) );
  COND1XL U16489 ( .A(n11978), .B(n16694), .C(n16686), .Z(n10153) );
  CANR2X1 U16490 ( .A(n16694), .B(poly14_shifted[270]), .C(n17598), .D(
        poly14_shifted[254]), .Z(n16687) );
  COND1XL U16491 ( .A(n13418), .B(n16694), .C(n16687), .Z(n10151) );
  CANR2X1 U16492 ( .A(n16694), .B(poly14_shifted[253]), .C(n17755), .D(
        poly14_shifted[237]), .Z(n16688) );
  COND1XL U16493 ( .A(n17065), .B(n16694), .C(n16688), .Z(n10168) );
  CANR2X1 U16494 ( .A(n16694), .B(poly14_shifted[251]), .C(n17174), .D(
        poly14_shifted[235]), .Z(n16689) );
  COND1XL U16495 ( .A(n16994), .B(n16694), .C(n16689), .Z(n10170) );
  CANR2XL U16496 ( .A(n16694), .B(poly14_shifted[260]), .C(n18017), .D(
        poly14_shifted[244]), .Z(n16690) );
  COND1XL U16497 ( .A(n17707), .B(n16694), .C(n16690), .Z(n10161) );
  CANR2X1 U16498 ( .A(n16694), .B(poly14_shifted[252]), .C(n16919), .D(
        poly14_shifted[236]), .Z(n16691) );
  COND1XL U16499 ( .A(n17087), .B(n16694), .C(n16691), .Z(n10169) );
  CANR2X1 U16500 ( .A(n16694), .B(poly14_shifted[254]), .C(n17099), .D(
        poly14_shifted[238]), .Z(n16692) );
  COND1XL U16501 ( .A(n12764), .B(n16694), .C(n16692), .Z(n10167) );
  CANR2X1 U16502 ( .A(n16694), .B(poly14_shifted[265]), .C(n16695), .D(
        poly14_shifted[249]), .Z(n16693) );
  COND1XL U16503 ( .A(n17123), .B(n16694), .C(n16693), .Z(n10156) );
  CANR2X1 U16504 ( .A(n16694), .B(poly14_shifted[249]), .C(n16695), .D(
        poly14_shifted[233]), .Z(n16696) );
  COND1XL U16505 ( .A(n17208), .B(n16694), .C(n16696), .Z(n10172) );
  CANR2X1 U16506 ( .A(n17990), .B(poly13_shifted[483]), .C(n18234), .D(
        poly13_shifted[469]), .Z(n16697) );
  COND1XL U16507 ( .A(n12006), .B(n17990), .C(n16697), .Z(n10591) );
  CANR2X1 U16508 ( .A(n17990), .B(poly13_shifted[465]), .C(poly13_shifted[451]), .D(n17755), .Z(n16698) );
  COND1XL U16509 ( .A(n13275), .B(n17990), .C(n16698), .Z(n10609) );
  CANR2X1 U16510 ( .A(n17990), .B(poly13_shifted[491]), .C(n17203), .D(
        poly13_shifted[477]), .Z(n16699) );
  COND1XL U16511 ( .A(n17185), .B(n17990), .C(n16699), .Z(n10583) );
  CANR2X1 U16512 ( .A(n17595), .B(poly13_shifted[249]), .C(n16700), .D(
        poly13_shifted[235]), .Z(n16701) );
  COND1XL U16513 ( .A(n16994), .B(n17595), .C(n16701), .Z(n10825) );
  CANR2X1 U16514 ( .A(n17990), .B(poly13_shifted[478]), .C(n16702), .D(
        poly13_shifted[464]), .Z(n16703) );
  COND1XL U16515 ( .A(n17062), .B(n17990), .C(n16703), .Z(n10596) );
  CANR2X1 U16516 ( .A(n17595), .B(poly13_shifted[244]), .C(n16326), .D(
        poly13_shifted[230]), .Z(n16704) );
  COND1XL U16517 ( .A(n16779), .B(n17595), .C(n16704), .Z(n10830) );
  CANR2X1 U16518 ( .A(n17595), .B(poly13_shifted[251]), .C(n17965), .D(
        poly13_shifted[237]), .Z(n16705) );
  COND1XL U16519 ( .A(n17065), .B(n17595), .C(n16705), .Z(n10823) );
  CANR2X1 U16520 ( .A(n17595), .B(poly13_shifted[247]), .C(n17755), .D(
        poly13_shifted[233]), .Z(n16706) );
  COND1XL U16521 ( .A(n17208), .B(n17595), .C(n16706), .Z(n10827) );
  CANR2X1 U16522 ( .A(n12185), .B(Poly11[25]), .C(n16644), .D(
        poly11_shifted[25]), .Z(n16707) );
  COND1XL U16523 ( .A(n17200), .B(n12185), .C(n16707), .Z(n11164) );
  CANR2X1 U16524 ( .A(n12185), .B(Poly11[21]), .C(n17533), .D(
        poly11_shifted[21]), .Z(n16708) );
  COND1XL U16525 ( .A(n17036), .B(n12185), .C(n16708), .Z(n11168) );
  CANR2X1 U16526 ( .A(n17755), .B(poly0_shifted[157]), .C(Poly0[157]), .D(
        n17671), .Z(n16709) );
  COND1XL U16527 ( .A(n17674), .B(n17185), .C(n16709), .Z(n9420) );
  CANR2X1 U16528 ( .A(n16644), .B(poly0_shifted[145]), .C(poly0_shifted[163]), 
        .D(n17671), .Z(n16710) );
  COND1XL U16529 ( .A(n17674), .B(n17076), .C(n16710), .Z(n9432) );
  CEOXL U16530 ( .A(Poly9[22]), .B(Poly9[111]), .Z(n16711) );
  CENX1 U16531 ( .A(Poly9[114]), .B(n16711), .Z(n16712) );
  CNR2XL U16532 ( .A(n17744), .B(n16712), .Z(n16713) );
  CANR1XL U16533 ( .A(poly9_shifted[44]), .B(n13351), .C(n16713), .Z(n16714)
         );
  COND1XL U16534 ( .A(n17711), .B(n13351), .C(n16714), .Z(n11272) );
  CANR2X1 U16535 ( .A(n17043), .B(Poly13[389]), .C(n17755), .D(
        poly13_shifted[389]), .Z(n16715) );
  COND1XL U16536 ( .A(n11995), .B(n17043), .C(n16715), .Z(n10671) );
  CANR2X1 U16537 ( .A(n17043), .B(Poly13[387]), .C(n17705), .D(
        poly13_shifted[387]), .Z(n16716) );
  COND1XL U16538 ( .A(n13275), .B(n17043), .C(n16716), .Z(n10673) );
  CEOXL U16539 ( .A(Poly13[526]), .B(Poly13[399]), .Z(n16717) );
  CANR2X1 U16540 ( .A(n17043), .B(poly13_shifted[427]), .C(n17755), .D(n16717), 
        .Z(n16718) );
  COND1XL U16541 ( .A(n17185), .B(n17043), .C(n16718), .Z(n10647) );
  CANR2X1 U16542 ( .A(n17043), .B(poly13_shifted[398]), .C(n17538), .D(
        poly13_shifted[384]), .Z(n16719) );
  COND1XL U16543 ( .A(n17751), .B(n17043), .C(n16719), .Z(n10676) );
  CANR2X1 U16544 ( .A(n16854), .B(poly8_shifted[75]), .C(poly12_shifted[124]), 
        .D(n16837), .Z(n16723) );
  CANR2X1 U16545 ( .A(n16867), .B(Poly4[44]), .C(n16874), .D(poly9_shifted[44]), .Z(n16722) );
  CANR2X1 U16546 ( .A(n16841), .B(poly8_shifted[68]), .C(n16866), .D(Poly5[80]), .Z(n16721) );
  CANR2X1 U16547 ( .A(n16840), .B(Poly6[16]), .C(n16862), .D(poly2_shifted[28]), .Z(n16720) );
  CANR2X1 U16548 ( .A(n16876), .B(poly5_shifted[38]), .C(n16839), .D(
        Poly15[32]), .Z(n16727) );
  CANR2X1 U16549 ( .A(n16875), .B(Poly2[38]), .C(n16855), .D(
        poly13_shifted[352]), .Z(n16726) );
  CANR2X1 U16550 ( .A(n16850), .B(Poly4[16]), .C(n16863), .D(Poly6[42]), .Z(
        n16725) );
  CANR2X1 U16551 ( .A(n16844), .B(Poly2[50]), .C(n16853), .D(
        poly13_shifted[390]), .Z(n16724) );
  CAN4X1 U16552 ( .A(n16727), .B(n16726), .C(n16725), .D(n16724), .Z(n16738)
         );
  CANR2X1 U16553 ( .A(n16838), .B(poly10_shifted[20]), .C(n12084), .D(
        Poly12[115]), .Z(n16731) );
  CIVXL U16554 ( .A(n16728), .Z(n16729) );
  CANR2X1 U16555 ( .A(n16842), .B(Poly3[39]), .C(Poly12[17]), .D(n16849), .Z(
        n16730) );
  CANR2X1 U16556 ( .A(n12071), .B(Poly14[285]), .C(n16865), .D(Poly11[83]), 
        .Z(n16735) );
  CANR2X1 U16557 ( .A(n16873), .B(Poly9[23]), .C(n16860), .D(poly5_shifted[57]), .Z(n16734) );
  CANR2X1 U16558 ( .A(n12067), .B(poly14_shifted[51]), .C(n16851), .D(
        Poly15[27]), .Z(n16733) );
  CANR2X1 U16559 ( .A(n16861), .B(poly8_shifted[58]), .C(n16877), .D(
        poly13_shifted[425]), .Z(n16732) );
  CAN4X1 U16560 ( .A(n16735), .B(n16734), .C(n16733), .D(n16732), .Z(n16736)
         );
  CIVXL U16561 ( .A(poly15_shifted[51]), .Z(n16745) );
  CEOXL U16562 ( .A(Poly15[47]), .B(Poly15[21]), .Z(n16739) );
  CEOXL U16563 ( .A(Poly15[53]), .B(n16739), .Z(n16743) );
  CANR11X1 U16564 ( .A(n18234), .B(n16743), .C(n16742), .D(n16741), .Z(n16744)
         );
  CANR2X1 U16565 ( .A(n16839), .B(Poly10[4]), .C(poly9_shifted[71]), .D(n16837), .Z(n16749) );
  CANR2X1 U16566 ( .A(n12071), .B(poly6_shifted[55]), .C(n16855), .D(
        Poly11[28]), .Z(n16748) );
  CANR2X1 U16567 ( .A(n16842), .B(poly13_shifted[507]), .C(n16872), .D(
        Poly11[73]), .Z(n16747) );
  CANR2X1 U16568 ( .A(n16849), .B(Poly10[20]), .C(n16852), .D(Poly11[63]), .Z(
        n16746) );
  CAN4X1 U16569 ( .A(n16749), .B(n16748), .C(n16747), .D(n16746), .Z(n16766)
         );
  CANR2X1 U16570 ( .A(n16838), .B(Poly4[20]), .C(n16851), .D(
        poly0_shifted[119]), .Z(n16752) );
  CANR2X1 U16571 ( .A(n12067), .B(poly5_shifted[88]), .C(n16841), .D(Poly2[30]), .Z(n16751) );
  CANR2X1 U16572 ( .A(n16875), .B(poly12_shifted[58]), .C(n16873), .D(
        poly7_shifted[330]), .Z(n16758) );
  CANR2X1 U16573 ( .A(n16876), .B(poly11_shifted[24]), .C(n16862), .D(
        Poly3[42]), .Z(n16757) );
  CIVXL U16574 ( .A(n16753), .Z(n16754) );
  CANR2X1 U16575 ( .A(n16866), .B(Poly11[72]), .C(n16754), .D(n16877), .Z(
        n16756) );
  CANR2X1 U16576 ( .A(n16867), .B(Poly15[57]), .C(n16854), .D(
        poly2_shifted[23]), .Z(n16755) );
  CAN4X1 U16577 ( .A(n16758), .B(n16757), .C(n16756), .D(n16755), .Z(n16764)
         );
  CANR2X1 U16578 ( .A(n16864), .B(Poly5[79]), .C(n12084), .D(Poly11[40]), .Z(
        n16762) );
  CANR2X1 U16579 ( .A(n16865), .B(poly8_shifted[72]), .C(n16853), .D(Poly5[86]), .Z(n16761) );
  CANR2X1 U16580 ( .A(n16860), .B(Poly10[25]), .C(n16843), .D(n17925), .Z(
        n16760) );
  CANR2X1 U16581 ( .A(n16861), .B(poly13_shifted[110]), .C(n16874), .D(
        poly15_shifted[22]), .Z(n16759) );
  CAN4X1 U16582 ( .A(n16762), .B(n16761), .C(n16760), .D(n16759), .Z(n16763)
         );
  CND4X1 U16583 ( .A(n16766), .B(n16765), .C(n16764), .D(n16763), .Z(n16767)
         );
  CAOR2XL U16584 ( .A(polydata[11]), .B(n17959), .C(n16767), .D(n16886), .Z(
        n8695) );
  CANR2X1 U16585 ( .A(n17977), .B(poly13_shifted[148]), .C(n17755), .D(
        poly13_shifted[134]), .Z(n16768) );
  COND1XL U16586 ( .A(n16779), .B(n17977), .C(n16768), .Z(n10926) );
  CANR2X1 U16587 ( .A(n17977), .B(poly13_shifted[158]), .C(n17523), .D(
        poly13_shifted[144]), .Z(n16769) );
  COND1XL U16588 ( .A(n17211), .B(n17977), .C(n16769), .Z(n10916) );
  CANR2X1 U16589 ( .A(n17977), .B(poly13_shifted[156]), .C(n17174), .D(
        poly13_shifted[142]), .Z(n16770) );
  COND1XL U16590 ( .A(n17699), .B(n17977), .C(n16770), .Z(n10918) );
  CANR2X1 U16591 ( .A(n17977), .B(Poly13[159]), .C(n17655), .D(
        poly13_shifted[159]), .Z(n16771) );
  COND1XL U16592 ( .A(n17188), .B(n17977), .C(n16771), .Z(n10901) );
  CANR2X1 U16593 ( .A(n17977), .B(poly13_shifted[145]), .C(n18047), .D(
        poly13_shifted[131]), .Z(n16772) );
  COND1XL U16594 ( .A(n13275), .B(n17977), .C(n16772), .Z(n10929) );
  CANR2X1 U16595 ( .A(n17977), .B(poly13_shifted[159]), .C(n17094), .D(
        poly13_shifted[145]), .Z(n16773) );
  COND1XL U16596 ( .A(n17173), .B(n17977), .C(n16773), .Z(n10915) );
  CANR2X1 U16597 ( .A(n17977), .B(poly13_shifted[144]), .C(n16919), .D(
        poly13_shifted[130]), .Z(n16774) );
  COND1XL U16598 ( .A(n16775), .B(n17977), .C(n16774), .Z(n10930) );
  CANR2X1 U16599 ( .A(n12958), .B(poly14_shifted[101]), .C(n17620), .D(
        poly14_shifted[85]), .Z(n16776) );
  COND1XL U16600 ( .A(n12006), .B(n12958), .C(n16776), .Z(n10320) );
  CANR2X1 U16601 ( .A(n12958), .B(poly14_shifted[90]), .C(n18234), .D(
        poly14_shifted[74]), .Z(n16777) );
  COND1XL U16602 ( .A(n12014), .B(n12958), .C(n16777), .Z(n10331) );
  CANR2X1 U16603 ( .A(n12958), .B(poly14_shifted[86]), .C(n17714), .D(
        poly14_shifted[70]), .Z(n16778) );
  COND1XL U16604 ( .A(n16779), .B(n12958), .C(n16778), .Z(n10335) );
  CANR2X1 U16605 ( .A(n12958), .B(poly14_shifted[100]), .C(n17705), .D(
        poly14_shifted[84]), .Z(n16780) );
  COND1XL U16606 ( .A(n16391), .B(n12958), .C(n16780), .Z(n10321) );
  CANR2X1 U16607 ( .A(n12958), .B(poly14_shifted[105]), .C(n17362), .D(
        poly14_shifted[89]), .Z(n16781) );
  COND1XL U16608 ( .A(n17123), .B(n12958), .C(n16781), .Z(n10316) );
  CANR2X1 U16609 ( .A(n12958), .B(poly14_shifted[92]), .C(n17504), .D(
        poly14_shifted[76]), .Z(n16782) );
  COND1XL U16610 ( .A(n17087), .B(n12958), .C(n16782), .Z(n10329) );
  CANR2X1 U16611 ( .A(n12958), .B(poly14_shifted[108]), .C(n17362), .D(
        poly14_shifted[92]), .Z(n16783) );
  COND1XL U16612 ( .A(n11978), .B(n12958), .C(n16783), .Z(n10313) );
  CANR2X1 U16613 ( .A(n12958), .B(poly14_shifted[102]), .C(n17714), .D(
        poly14_shifted[86]), .Z(n16784) );
  COND1XL U16614 ( .A(n17753), .B(n12958), .C(n16784), .Z(n10319) );
  CANR2X1 U16615 ( .A(n12958), .B(poly14_shifted[95]), .C(n17965), .D(
        poly14_shifted[79]), .Z(n16785) );
  COND1XL U16616 ( .A(n17196), .B(n12958), .C(n16785), .Z(n10326) );
  CANR2X1 U16617 ( .A(n12958), .B(poly14_shifted[111]), .C(n17535), .D(
        poly14_shifted[95]), .Z(n16786) );
  COND1XL U16618 ( .A(n17188), .B(n12958), .C(n16786), .Z(n10310) );
  CANR2X1 U16619 ( .A(n12958), .B(poly14_shifted[88]), .C(n16787), .D(
        poly14_shifted[72]), .Z(n16788) );
  COND1XL U16620 ( .A(n17166), .B(n12958), .C(n16788), .Z(n10333) );
  CANR2X1 U16621 ( .A(n17332), .B(Poly1[336]), .C(n18047), .D(
        poly1_shifted[336]), .Z(n16789) );
  COND1XL U16622 ( .A(n17062), .B(n17332), .C(n16789), .Z(n9021) );
  CANR2X1 U16623 ( .A(n17332), .B(Poly1[337]), .C(n17560), .D(
        poly1_shifted[337]), .Z(n16790) );
  COND1XL U16624 ( .A(n17173), .B(n17332), .C(n16790), .Z(n9020) );
  CANR2X1 U16625 ( .A(n17332), .B(Poly1[340]), .C(n17560), .D(
        poly1_shifted[340]), .Z(n16791) );
  COND1XL U16626 ( .A(n16391), .B(n17332), .C(n16791), .Z(n9017) );
  CANR2X1 U16627 ( .A(n17332), .B(poly1_shifted[343]), .C(n18234), .D(
        poly1_shifted[332]), .Z(n16792) );
  COND1XL U16628 ( .A(n17087), .B(n17332), .C(n16792), .Z(n9025) );
  CANR2X1 U16629 ( .A(n18028), .B(poly7_shifted[330]), .C(n17545), .D(
        poly7_shifted[318]), .Z(n16793) );
  COND1XL U16630 ( .A(n13418), .B(n18028), .C(n16793), .Z(n9786) );
  CANR2X1 U16631 ( .A(n18028), .B(poly7_shifted[325]), .C(n17535), .D(
        poly7_shifted[313]), .Z(n16794) );
  COND1XL U16632 ( .A(n17200), .B(n18028), .C(n16794), .Z(n9791) );
  CANR2XL U16633 ( .A(n13351), .B(poly9_shifted[69]), .C(poly9_shifted[58]), 
        .D(n18017), .Z(n16795) );
  COND1XL U16634 ( .A(n17735), .B(n13351), .C(n16795), .Z(n11247) );
  CANR2X1 U16635 ( .A(n16873), .B(n18220), .C(n16796), .D(n16840), .Z(n16800)
         );
  CANR2X1 U16636 ( .A(n16861), .B(Poly6[29]), .C(n16874), .D(poly7_shifted[85]), .Z(n16799) );
  CANR2X1 U16637 ( .A(n16863), .B(poly1_shifted[114]), .C(n16852), .D(
        poly8_shifted[44]), .Z(n16798) );
  CANR2X1 U16638 ( .A(n16843), .B(Poly10[22]), .C(n16862), .D(
        poly5_shifted[34]), .Z(n16797) );
  CAN4X1 U16639 ( .A(n16800), .B(n16799), .C(n16798), .D(n16797), .Z(n16815)
         );
  CANR2X1 U16640 ( .A(n16876), .B(poly10_shifted[17]), .C(Poly15[33]), .D(
        n16837), .Z(n16805) );
  CANR2X1 U16641 ( .A(n16850), .B(Poly6[1]), .C(n16877), .D(Poly4[32]), .Z(
        n16804) );
  CANR2X1 U16642 ( .A(n12067), .B(Poly6[18]), .C(n16801), .D(n16838), .Z(
        n16803) );
  CANR2X1 U16643 ( .A(n16875), .B(Poly6[43]), .C(n16867), .D(
        poly14_shifted[66]), .Z(n16802) );
  CAN4X1 U16644 ( .A(n16805), .B(n16804), .C(n16803), .D(n16802), .Z(n16814)
         );
  CANR2X1 U16645 ( .A(n16842), .B(poly2_shifted[20]), .C(n16839), .D(
        poly0_shifted[218]), .Z(n16807) );
  CANR2X1 U16646 ( .A(n16865), .B(poly0_shifted[49]), .C(n16860), .D(Poly4[37]), .Z(n16806) );
  CANR2X1 U16647 ( .A(n12071), .B(poly7_shifted[59]), .C(n12084), .D(
        Poly15[13]), .Z(n16811) );
  CANR2X1 U16648 ( .A(n16853), .B(Poly4[34]), .C(n16851), .D(Poly9[89]), .Z(
        n16810) );
  CANR2X1 U16649 ( .A(n16844), .B(poly13_shifted[399]), .C(n16841), .D(
        Poly4[23]), .Z(n16809) );
  CANR2X1 U16650 ( .A(n16849), .B(Poly11[25]), .C(n16872), .D(
        poly4_shifted[31]), .Z(n16808) );
  CAN4X1 U16651 ( .A(n16811), .B(n16810), .C(n16809), .D(n16808), .Z(n16812)
         );
  CND4X1 U16652 ( .A(n16815), .B(n16814), .C(n16813), .D(n16812), .Z(n16816)
         );
  CAOR2XL U16653 ( .A(polydata[6]), .B(n17495), .C(n16816), .D(n16886), .Z(
        n8690) );
  CANR2X1 U16654 ( .A(n16850), .B(Poly10[31]), .C(n16873), .D(
        poly0_shifted[208]), .Z(n16821) );
  CANR2X1 U16655 ( .A(n12084), .B(poly0_shifted[52]), .C(n16872), .D(
        poly3_shifted[39]), .Z(n16820) );
  CANR2X1 U16656 ( .A(n16876), .B(poly1_shifted[96]), .C(n16851), .D(
        poly4_shifted[28]), .Z(n16819) );
  CIVX1 U16657 ( .A(n16817), .Z(n17957) );
  CANR2X1 U16658 ( .A(n16864), .B(n17957), .C(poly1_shifted[127]), .D(n16862), 
        .Z(n16818) );
  CAN4X1 U16659 ( .A(n16821), .B(n16820), .C(n16819), .D(n16818), .Z(n16835)
         );
  CANR2X1 U16660 ( .A(n16844), .B(Poly11[81]), .C(n16843), .D(Poly3[41]), .Z(
        n16825) );
  CANR2X1 U16661 ( .A(n16842), .B(poly1_shifted[233]), .C(n16860), .D(
        Poly2[58]), .Z(n16824) );
  CANR2X1 U16662 ( .A(n16854), .B(Poly6[19]), .C(n16877), .D(Poly12[29]), .Z(
        n16823) );
  CANR2X1 U16663 ( .A(n16840), .B(Poly11[74]), .C(poly1_shifted[131]), .D(
        n16849), .Z(n16822) );
  CAN4X1 U16664 ( .A(n16825), .B(n16824), .C(n16823), .D(n16822), .Z(n16834)
         );
  CANR2X1 U16665 ( .A(n16852), .B(poly7_shifted[159]), .C(Poly4[45]), .D(
        n16837), .Z(n16829) );
  CANR2X1 U16666 ( .A(n16838), .B(Poly11[68]), .C(n16874), .D(Poly2[25]), .Z(
        n16828) );
  CANR2X1 U16667 ( .A(n16863), .B(Poly13[394]), .C(n16866), .D(Poly3[81]), .Z(
        n16827) );
  CANR2X1 U16668 ( .A(n16861), .B(poly3_shifted[36]), .C(n16867), .D(
        poly5_shifted[40]), .Z(n16826) );
  CAN4X1 U16669 ( .A(n16829), .B(n16828), .C(n16827), .D(n16826), .Z(n16833)
         );
  CANR2X1 U16670 ( .A(n12071), .B(poly1_shifted[47]), .C(n16839), .D(
        poly12_shifted[89]), .Z(n16831) );
  CANR2X1 U16671 ( .A(n16865), .B(Poly6[4]), .C(n16841), .D(
        poly14_shifted[297]), .Z(n16830) );
  CND4X1 U16672 ( .A(n16835), .B(n16834), .C(n16833), .D(n16832), .Z(n16836)
         );
  CAOR2XL U16673 ( .A(polydata[7]), .B(n17959), .C(n16836), .D(n16886), .Z(
        n8691) );
  CANR2X1 U16674 ( .A(n16838), .B(poly7_shifted[164]), .C(poly8_shifted[73]), 
        .D(n16837), .Z(n16848) );
  CANR2X1 U16675 ( .A(n16840), .B(Poly12[31]), .C(n16839), .D(Poly4[38]), .Z(
        n16847) );
  CANR2X1 U16676 ( .A(n16842), .B(poly14_shifted[170]), .C(n16841), .D(
        Poly10[12]), .Z(n16846) );
  CANR2X1 U16677 ( .A(n16844), .B(poly9_shifted[55]), .C(n16843), .D(
        poly0_shifted[217]), .Z(n16845) );
  CAN4X1 U16678 ( .A(n16848), .B(n16847), .C(n16846), .D(n16845), .Z(n16885)
         );
  CANR2X1 U16679 ( .A(n16850), .B(poly8_shifted[32]), .C(poly5_shifted[49]), 
        .D(n16849), .Z(n16859) );
  CANR2X1 U16680 ( .A(n12084), .B(poly9_shifted[76]), .C(n16851), .D(Poly6[25]), .Z(n16858) );
  CANR2X1 U16681 ( .A(n16853), .B(poly14_shifted[155]), .C(n16852), .D(
        Poly12[58]), .Z(n16857) );
  CANR2X1 U16682 ( .A(n16855), .B(Poly1[61]), .C(n16854), .D(Poly0[211]), .Z(
        n16856) );
  CAN4X1 U16683 ( .A(n16859), .B(n16858), .C(n16857), .D(n16856), .Z(n16884)
         );
  CANR2X1 U16684 ( .A(n16861), .B(poly5_shifted[22]), .C(n16860), .D(
        Poly15[12]), .Z(n16871) );
  CANR2X1 U16685 ( .A(n16863), .B(poly7_shifted[332]), .C(n16862), .D(
        Poly4[30]), .Z(n16870) );
  CANR2X2 U16686 ( .A(n16865), .B(Poly14[205]), .C(n16864), .D(
        poly15_shifted[50]), .Z(n16869) );
  CANR2X1 U16687 ( .A(n16867), .B(poly9_shifted[87]), .C(n16866), .D(
        poly2_shifted[13]), .Z(n16868) );
  CAN4X1 U16688 ( .A(n16871), .B(n16870), .C(n16869), .D(n16868), .Z(n16883)
         );
  CANR2X1 U16689 ( .A(n16873), .B(poly14_shifted[78]), .C(n16872), .D(
        Poly15[16]), .Z(n16881) );
  CANR2X1 U16690 ( .A(n16875), .B(poly8_shifted[66]), .C(n16874), .D(
        Poly12[91]), .Z(n16880) );
  CANR2X1 U16691 ( .A(n12071), .B(poly9_shifted[42]), .C(n16876), .D(
        poly9_shifted[111]), .Z(n16879) );
  CANR2X1 U16692 ( .A(n12067), .B(poly1_shifted[265]), .C(n16877), .D(
        Poly6[14]), .Z(n16878) );
  CAN4X1 U16693 ( .A(n16881), .B(n16880), .C(n16879), .D(n16878), .Z(n16882)
         );
  CND4X1 U16694 ( .A(n16885), .B(n16884), .C(n16883), .D(n16882), .Z(n16887)
         );
  CAOR2XL U16695 ( .A(polydata[8]), .B(n17495), .C(n16887), .D(n16886), .Z(
        n8692) );
  CANR2X1 U16696 ( .A(n18044), .B(Poly15[20]), .C(n17655), .D(
        poly15_shifted[20]), .Z(n16888) );
  COND1XL U16697 ( .A(n17707), .B(n18044), .C(n16888), .Z(n9617) );
  CANR2X1 U16698 ( .A(n18044), .B(Poly15[17]), .C(n17375), .D(
        poly15_shifted[17]), .Z(n16889) );
  COND1XL U16699 ( .A(n17173), .B(n18044), .C(n16889), .Z(n9620) );
  CANR2X1 U16700 ( .A(n18044), .B(poly15_shifted[22]), .C(n17094), .D(
        Poly15[52]), .Z(n16890) );
  COND1XL U16701 ( .A(n16939), .B(n18044), .C(n16890), .Z(n9630) );
  CANR2X1 U16702 ( .A(n18044), .B(Poly15[12]), .C(n17352), .D(Poly15[57]), .Z(
        n16891) );
  COND1XL U16703 ( .A(n17087), .B(n18044), .C(n16891), .Z(n9625) );
  CANR2X1 U16704 ( .A(n18044), .B(poly15_shifted[25]), .C(n16326), .D(
        Poly15[55]), .Z(n16892) );
  COND1XL U16705 ( .A(n12014), .B(n18044), .C(n16892), .Z(n9627) );
  CANR2X1 U16706 ( .A(n18044), .B(poly15_shifted[15]), .C(n17613), .D(
        Poly15[45]), .Z(n16893) );
  COND1XL U16707 ( .A(n17751), .B(n18044), .C(n16893), .Z(n9637) );
  CANR2X1 U16708 ( .A(n18044), .B(Poly15[24]), .C(n17198), .D(
        poly15_shifted[24]), .Z(n16894) );
  COND1XL U16709 ( .A(n17721), .B(n18044), .C(n16894), .Z(n9613) );
  CANR2X1 U16710 ( .A(n18044), .B(poly15_shifted[26]), .C(n16435), .D(
        Poly15[56]), .Z(n16895) );
  COND1XL U16711 ( .A(n16994), .B(n18044), .C(n16895), .Z(n9626) );
  CANR2X1 U16712 ( .A(n18044), .B(Poly15[16]), .C(n17527), .D(
        poly15_shifted[16]), .Z(n16896) );
  COND1XL U16713 ( .A(n17211), .B(n18044), .C(n16896), .Z(n9621) );
  CANR2X1 U16714 ( .A(n18044), .B(poly15_shifted[21]), .C(n17375), .D(
        Poly15[51]), .Z(n16897) );
  COND1XL U16715 ( .A(n17757), .B(n18044), .C(n16897), .Z(n9631) );
  CANR2X1 U16716 ( .A(n18044), .B(poly15_shifted[20]), .C(n17198), .D(
        Poly15[50]), .Z(n16898) );
  COND1XL U16717 ( .A(n11995), .B(n18044), .C(n16898), .Z(n9632) );
  CANR2X1 U16718 ( .A(n18044), .B(Poly15[21]), .C(n17375), .D(
        poly15_shifted[21]), .Z(n16899) );
  COND1XL U16719 ( .A(n12006), .B(n18044), .C(n16899), .Z(n9616) );
  CANR2X1 U16720 ( .A(n18044), .B(poly15_shifted[23]), .C(n17352), .D(
        Poly15[53]), .Z(n16900) );
  COND1XL U16721 ( .A(n17163), .B(n18044), .C(n16900), .Z(n9629) );
  CEOXL U16722 ( .A(Poly15[12]), .B(Poly15[45]), .Z(n16901) );
  CANR2X1 U16723 ( .A(n18044), .B(Poly15[27]), .C(n17352), .D(n16901), .Z(
        n16902) );
  COND1XL U16724 ( .A(n17741), .B(n18044), .C(n16902), .Z(n9610) );
  CANR2X1 U16725 ( .A(n13070), .B(poly7_shifted[159]), .C(n17552), .D(
        poly7_shifted[147]), .Z(n16903) );
  COND1XL U16726 ( .A(n17658), .B(n13070), .C(n16903), .Z(n9957) );
  CANR2X1 U16727 ( .A(n17072), .B(poly0_shifted[155]), .C(n17671), .D(
        Poly0[155]), .Z(n16904) );
  COND1XL U16728 ( .A(n17674), .B(n17741), .C(n16904), .Z(n9422) );
  CANR2X1 U16729 ( .A(n17755), .B(poly0_shifted[158]), .C(n17671), .D(
        Poly0[158]), .Z(n16905) );
  COND1XL U16730 ( .A(n17674), .B(n17004), .C(n16905), .Z(n9419) );
  CEOX1 U16731 ( .A(n16907), .B(n16906), .Z(n16908) );
  CENX1 U16732 ( .A(Poly4[28]), .B(n16908), .Z(n16910) );
  CMXI2XL U16733 ( .A0(n18219), .A1(Poly4[45]), .S(n12153), .Z(n16909) );
  COND1XL U16734 ( .A(n16910), .B(n17744), .C(n16909), .Z(n8811) );
  CANR2X1 U16735 ( .A(n16985), .B(poly3_shifted[80]), .C(Poly3[80]), .D(n17359), .Z(n16911) );
  COND1XL U16736 ( .A(n17361), .B(n17062), .C(n16911), .Z(n8860) );
  CANR2X1 U16737 ( .A(n17714), .B(poly3_shifted[81]), .C(Poly3[81]), .D(n17359), .Z(n16912) );
  COND1XL U16738 ( .A(n17361), .B(n17076), .C(n16912), .Z(n8859) );
  CANR2X1 U16739 ( .A(n17714), .B(poly3_shifted[76]), .C(Poly3[76]), .D(n17359), .Z(n16913) );
  COND1XL U16740 ( .A(n17361), .B(n17087), .C(n16913), .Z(n8864) );
  CANR2XL U16741 ( .A(n17755), .B(poly3_shifted[74]), .C(Poly3[74]), .D(n17359), .Z(n16914) );
  COND1XL U16742 ( .A(n17361), .B(n12014), .C(n16914), .Z(n8866) );
  CANR2X1 U16743 ( .A(n17508), .B(poly3_shifted[73]), .C(Poly3[73]), .D(n17359), .Z(n16915) );
  COND1XL U16744 ( .A(n17361), .B(n17208), .C(n16915), .Z(n8867) );
  CANR2X1 U16745 ( .A(n13351), .B(poly9_shifted[58]), .C(n17238), .D(
        poly9_shifted[47]), .Z(n16916) );
  COND1XL U16746 ( .A(n17196), .B(n13351), .C(n16916), .Z(n11258) );
  CANR2X1 U16747 ( .A(n13351), .B(poly9_shifted[73]), .C(n17072), .D(
        poly9_shifted[62]), .Z(n16917) );
  COND1XL U16748 ( .A(n13418), .B(n13351), .C(n16917), .Z(n11243) );
  CANR2X1 U16749 ( .A(n16787), .B(poly0_shifted[148]), .C(n17671), .D(
        poly0_shifted[166]), .Z(n16918) );
  COND1XL U16750 ( .A(n17674), .B(n16391), .C(n16918), .Z(n9429) );
  CANR2X1 U16751 ( .A(n16919), .B(poly0_shifted[143]), .C(n17671), .D(
        poly0_shifted[161]), .Z(n16920) );
  COND1XL U16752 ( .A(n17674), .B(n17196), .C(n16920), .Z(n9434) );
  CANR2X1 U16753 ( .A(n17504), .B(poly0_shifted[140]), .C(n17671), .D(
        poly0_shifted[158]), .Z(n16921) );
  COND1XL U16754 ( .A(n17674), .B(n17087), .C(n16921), .Z(n9437) );
  CANR2X1 U16755 ( .A(n17072), .B(poly0_shifted[159]), .C(n17671), .D(
        Poly0[159]), .Z(n16922) );
  COND1XL U16756 ( .A(n17674), .B(n17188), .C(n16922), .Z(n9418) );
  CANR2X1 U16757 ( .A(n17266), .B(poly0_shifted[144]), .C(n17671), .D(
        poly0_shifted[162]), .Z(n16923) );
  COND1XL U16758 ( .A(n17674), .B(n17062), .C(n16923), .Z(n9433) );
  CANR2X1 U16759 ( .A(n12977), .B(poly7_shifted[183]), .C(n17458), .D(
        poly7_shifted[171]), .Z(n16924) );
  COND1XL U16760 ( .A(n16994), .B(n12977), .C(n16924), .Z(n9933) );
  CANR2X1 U16761 ( .A(n12977), .B(poly7_shifted[187]), .C(n18234), .D(
        poly7_shifted[175]), .Z(n16925) );
  COND1XL U16762 ( .A(n17196), .B(n12977), .C(n16925), .Z(n9929) );
  CANR2X1 U16763 ( .A(n12977), .B(Poly7[182]), .C(n17290), .D(
        poly7_shifted[182]), .Z(n16926) );
  COND1XL U16764 ( .A(n17753), .B(n12977), .C(n16926), .Z(n9922) );
  CANR2X1 U16765 ( .A(n12977), .B(poly7_shifted[174]), .C(n17288), .D(
        poly7_shifted[162]), .Z(n16927) );
  COND1XL U16766 ( .A(n16775), .B(n12977), .C(n16927), .Z(n9942) );
  CANR2X1 U16767 ( .A(n12977), .B(poly7_shifted[175]), .C(n18234), .D(
        poly7_shifted[163]), .Z(n16928) );
  COND1XL U16768 ( .A(n13275), .B(n12977), .C(n16928), .Z(n9941) );
  CANR2X1 U16769 ( .A(n12977), .B(Poly7[187]), .C(n17598), .D(
        poly7_shifted[187]), .Z(n16929) );
  COND1XL U16770 ( .A(n17741), .B(n12977), .C(n16929), .Z(n9917) );
  CANR2X1 U16771 ( .A(n12977), .B(poly7_shifted[186]), .C(n17288), .D(
        poly7_shifted[174]), .Z(n16930) );
  COND1XL U16772 ( .A(n12764), .B(n12977), .C(n16930), .Z(n9930) );
  CANR2X1 U16773 ( .A(n12977), .B(Poly7[181]), .C(n17178), .D(
        poly7_shifted[181]), .Z(n16931) );
  COND1XL U16774 ( .A(n12006), .B(n12977), .C(n16931), .Z(n9923) );
  CANR2X1 U16775 ( .A(n12977), .B(Poly7[189]), .C(n17203), .D(
        poly7_shifted[189]), .Z(n16932) );
  COND1XL U16776 ( .A(n17185), .B(n12977), .C(n16932), .Z(n9915) );
  CANR2X1 U16777 ( .A(n17982), .B(poly13_shifted[373]), .C(poly13_shifted[359]), .D(n16947), .Z(n16933) );
  COND1XL U16778 ( .A(n17718), .B(n17982), .C(n16933), .Z(n10701) );
  CANR2X1 U16779 ( .A(n17603), .B(poly13_shifted[342]), .C(n17538), .D(
        poly13_shifted[328]), .Z(n16934) );
  COND1XL U16780 ( .A(n17166), .B(n17603), .C(n16934), .Z(n10732) );
  CANR2X1 U16781 ( .A(n17603), .B(poly13_shifted[355]), .C(n17298), .D(
        poly13_shifted[341]), .Z(n16935) );
  COND1XL U16782 ( .A(n12006), .B(n17603), .C(n16935), .Z(n10719) );
  CANR2X1 U16783 ( .A(n17603), .B(poly13_shifted[356]), .C(n17538), .D(
        poly13_shifted[342]), .Z(n16936) );
  COND1XL U16784 ( .A(n17001), .B(n17603), .C(n16936), .Z(n10718) );
  CANR2X1 U16785 ( .A(n17603), .B(poly13_shifted[343]), .C(n17298), .D(
        poly13_shifted[329]), .Z(n16937) );
  COND1XL U16786 ( .A(n17208), .B(n17603), .C(n16937), .Z(n10731) );
  CANR2X1 U16787 ( .A(n17603), .B(poly13_shifted[341]), .C(n17298), .D(
        poly13_shifted[327]), .Z(n16938) );
  COND1XL U16788 ( .A(n16939), .B(n17603), .C(n16938), .Z(n10733) );
  CANR2X1 U16789 ( .A(n17603), .B(poly13_shifted[347]), .C(n17755), .D(
        poly13_shifted[333]), .Z(n16940) );
  COND1XL U16790 ( .A(n17065), .B(n17603), .C(n16940), .Z(n10727) );
  CANR2X1 U16791 ( .A(n17603), .B(poly13_shifted[336]), .C(n17640), .D(
        poly13_shifted[322]), .Z(n16941) );
  COND1XL U16792 ( .A(n16775), .B(n17603), .C(n16941), .Z(n10738) );
  CANR2X1 U16793 ( .A(n17603), .B(poly13_shifted[346]), .C(n17965), .D(
        poly13_shifted[332]), .Z(n16942) );
  COND1XL U16794 ( .A(n17218), .B(n17603), .C(n16942), .Z(n10728) );
  CANR2X1 U16795 ( .A(n17603), .B(poly13_shifted[361]), .C(n17755), .D(
        poly13_shifted[347]), .Z(n16943) );
  COND1XL U16796 ( .A(n17741), .B(n17603), .C(n16943), .Z(n10713) );
  CANR2X1 U16797 ( .A(n17603), .B(poly13_shifted[349]), .C(n17613), .D(
        poly13_shifted[335]), .Z(n16944) );
  COND1XL U16798 ( .A(n17196), .B(n17603), .C(n16944), .Z(n10725) );
  CANR2X1 U16799 ( .A(n17603), .B(poly13_shifted[344]), .C(n17538), .D(
        poly13_shifted[330]), .Z(n16945) );
  COND1XL U16800 ( .A(n12014), .B(n17603), .C(n16945), .Z(n10730) );
  CANR2X1 U16801 ( .A(n17603), .B(poly13_shifted[337]), .C(n16644), .D(
        poly13_shifted[323]), .Z(n16946) );
  COND1XL U16802 ( .A(n13275), .B(n17603), .C(n16946), .Z(n10737) );
  CANR2X1 U16803 ( .A(n17603), .B(poly13_shifted[359]), .C(poly13_shifted[345]), .D(n16947), .Z(n16948) );
  COND1XL U16804 ( .A(n17123), .B(n17603), .C(n16948), .Z(n10715) );
  CANR2X1 U16805 ( .A(n17603), .B(poly13_shifted[335]), .C(n17613), .D(
        poly13_shifted[321]), .Z(n16949) );
  COND1XL U16806 ( .A(n16950), .B(n17603), .C(n16949), .Z(n10739) );
  CANR2X1 U16807 ( .A(n17603), .B(poly13_shifted[362]), .C(n17755), .D(
        poly13_shifted[348]), .Z(n16951) );
  COND1XL U16808 ( .A(n11978), .B(n17603), .C(n16951), .Z(n10712) );
  CANR2X1 U16809 ( .A(n17603), .B(poly13_shifted[364]), .C(n17705), .D(
        poly13_shifted[350]), .Z(n16952) );
  COND1XL U16810 ( .A(n13418), .B(n17603), .C(n16952), .Z(n10710) );
  CANR2X1 U16811 ( .A(n17603), .B(poly13_shifted[334]), .C(n17634), .D(
        poly13_shifted[320]), .Z(n16953) );
  COND1XL U16812 ( .A(n12011), .B(n17603), .C(n16953), .Z(n10740) );
  CANR2X1 U16813 ( .A(n17603), .B(poly13_shifted[363]), .C(n17613), .D(
        poly13_shifted[349]), .Z(n16954) );
  COND1XL U16814 ( .A(n17185), .B(n17603), .C(n16954), .Z(n10711) );
  CANR2X1 U16815 ( .A(n17603), .B(poly13_shifted[348]), .C(n17755), .D(
        poly13_shifted[334]), .Z(n16955) );
  COND1XL U16816 ( .A(n12764), .B(n17603), .C(n16955), .Z(n10726) );
  CNR2X1 U16817 ( .A(Poly6[18]), .B(n16956), .Z(n16960) );
  CNR2XL U16818 ( .A(n16957), .B(n16960), .Z(n16958) );
  CANR2X1 U16819 ( .A(n12206), .B(poly7_shifted[364]), .C(n17965), .D(
        poly7_shifted[352]), .Z(n16963) );
  COND1XL U16820 ( .A(n12011), .B(n12206), .C(n16963), .Z(n9752) );
  CANR2X1 U16821 ( .A(n12206), .B(poly7_shifted[385]), .C(n17535), .D(
        poly7_shifted[373]), .Z(n16964) );
  COND1XL U16822 ( .A(n12006), .B(n12206), .C(n16964), .Z(n9731) );
  CANR2X1 U16823 ( .A(n12206), .B(poly7_shifted[374]), .C(n17466), .D(
        poly7_shifted[362]), .Z(n16965) );
  COND1XL U16824 ( .A(n12014), .B(n12206), .C(n16965), .Z(n9742) );
  CANR2X1 U16825 ( .A(n12206), .B(poly7_shifted[393]), .C(n17121), .D(
        poly7_shifted[381]), .Z(n16966) );
  COND1XL U16826 ( .A(n17185), .B(n12206), .C(n16966), .Z(n9723) );
  CANR2X1 U16827 ( .A(n12206), .B(poly7_shifted[375]), .C(n17398), .D(
        poly7_shifted[363]), .Z(n16967) );
  COND1XL U16828 ( .A(n16994), .B(n12206), .C(n16967), .Z(n9741) );
  CANR2X1 U16829 ( .A(n12206), .B(poly7_shifted[384]), .C(n17535), .D(
        poly7_shifted[372]), .Z(n16968) );
  COND1XL U16830 ( .A(n16391), .B(n12206), .C(n16968), .Z(n9732) );
  CANR2X1 U16831 ( .A(n12206), .B(poly7_shifted[395]), .C(n17458), .D(
        poly7_shifted[383]), .Z(n16969) );
  COND1XL U16832 ( .A(n17188), .B(n12206), .C(n16969), .Z(n9721) );
  CANR2X1 U16833 ( .A(n12206), .B(poly7_shifted[372]), .C(n17535), .D(
        poly7_shifted[360]), .Z(n16970) );
  COND1XL U16834 ( .A(n17166), .B(n12206), .C(n16970), .Z(n9744) );
  CANR2X1 U16835 ( .A(n12206), .B(poly7_shifted[369]), .C(n17121), .D(
        poly7_shifted[357]), .Z(n16971) );
  COND1XL U16836 ( .A(n11993), .B(n12206), .C(n16971), .Z(n9747) );
  CANR2X1 U16837 ( .A(n12206), .B(poly7_shifted[367]), .C(n17453), .D(
        poly7_shifted[355]), .Z(n16972) );
  COND1XL U16838 ( .A(n13275), .B(n12206), .C(n16972), .Z(n9749) );
  CANR2X1 U16839 ( .A(n12206), .B(poly7_shifted[381]), .C(n17121), .D(
        poly7_shifted[369]), .Z(n16973) );
  COND1XL U16840 ( .A(n17173), .B(n12206), .C(n16973), .Z(n9735) );
  CANR2X1 U16841 ( .A(n12206), .B(poly7_shifted[379]), .C(n17453), .D(
        poly7_shifted[367]), .Z(n16974) );
  COND1XL U16842 ( .A(n17196), .B(n12206), .C(n16974), .Z(n9737) );
  CANR2X1 U16843 ( .A(n12206), .B(poly7_shifted[380]), .C(n17390), .D(
        poly7_shifted[368]), .Z(n16975) );
  COND1XL U16844 ( .A(n17211), .B(n12206), .C(n16975), .Z(n9736) );
  CANR2X1 U16845 ( .A(n12206), .B(poly7_shifted[386]), .C(n18047), .D(
        poly7_shifted[374]), .Z(n16976) );
  COND1XL U16846 ( .A(n17753), .B(n12206), .C(n16976), .Z(n9730) );
  CANR2X1 U16847 ( .A(n12206), .B(poly7_shifted[377]), .C(n17174), .D(
        poly7_shifted[365]), .Z(n16977) );
  COND1XL U16848 ( .A(n17065), .B(n12206), .C(n16977), .Z(n9739) );
  CANR2X1 U16849 ( .A(n12206), .B(poly7_shifted[378]), .C(n16372), .D(
        poly7_shifted[366]), .Z(n16978) );
  COND1XL U16850 ( .A(n12764), .B(n12206), .C(n16978), .Z(n9738) );
  CANR2X1 U16851 ( .A(n12206), .B(poly7_shifted[394]), .C(n17105), .D(
        poly7_shifted[382]), .Z(n16979) );
  COND1XL U16852 ( .A(n13418), .B(n12206), .C(n16979), .Z(n9722) );
  CANR2X1 U16853 ( .A(n12206), .B(poly7_shifted[365]), .C(n17174), .D(
        poly7_shifted[353]), .Z(n16980) );
  COND1XL U16854 ( .A(n16950), .B(n12206), .C(n16980), .Z(n9751) );
  CANR2X1 U16855 ( .A(n12206), .B(poly7_shifted[366]), .C(n17449), .D(
        poly7_shifted[354]), .Z(n16981) );
  COND1XL U16856 ( .A(n16303), .B(n12206), .C(n16981), .Z(n9750) );
  CANR2X1 U16857 ( .A(n12206), .B(poly7_shifted[370]), .C(n16323), .D(
        poly7_shifted[358]), .Z(n16982) );
  COND1XL U16858 ( .A(n17757), .B(n12206), .C(n16982), .Z(n9746) );
  CANR2X1 U16859 ( .A(n12206), .B(poly7_shifted[392]), .C(n17390), .D(
        poly7_shifted[380]), .Z(n16983) );
  COND1XL U16860 ( .A(n11978), .B(n12206), .C(n16983), .Z(n9724) );
  CANR2X1 U16861 ( .A(n12206), .B(poly7_shifted[389]), .C(n17174), .D(
        poly7_shifted[377]), .Z(n16984) );
  COND1XL U16862 ( .A(n17123), .B(n12206), .C(n16984), .Z(n9727) );
  CANR2X1 U16863 ( .A(n12206), .B(poly7_shifted[376]), .C(n16985), .D(
        poly7_shifted[364]), .Z(n16986) );
  COND1XL U16864 ( .A(n17087), .B(n12206), .C(n16986), .Z(n9740) );
  CANR2X1 U16865 ( .A(n12206), .B(poly7_shifted[388]), .C(n17343), .D(
        poly7_shifted[376]), .Z(n16987) );
  COND1XL U16866 ( .A(n16179), .B(n12206), .C(n16987), .Z(n9728) );
  CIVXL U16867 ( .A(n16988), .Z(n16990) );
  CMXI2XL U16868 ( .A0(n12004), .A1(poly4_shifted[21]), .S(n18230), .Z(n16989)
         );
  COND1XL U16869 ( .A(n17959), .B(n16990), .C(n16989), .Z(n8852) );
  CANR2X1 U16870 ( .A(n17969), .B(poly13_shifted[79]), .C(n17668), .D(
        poly13_shifted[65]), .Z(n16991) );
  COND1XL U16871 ( .A(n17697), .B(n17969), .C(n16991), .Z(n10995) );
  CANR2X1 U16872 ( .A(n17969), .B(poly13_shifted[107]), .C(n17668), .D(
        poly13_shifted[93]), .Z(n16992) );
  COND1XL U16873 ( .A(n17185), .B(n17969), .C(n16992), .Z(n10967) );
  CANR2X1 U16874 ( .A(n17620), .B(Poly0[213]), .C(Poly0[11]), .D(n17503), .Z(
        n16993) );
  COND1XL U16875 ( .A(n17506), .B(n16994), .C(n16993), .Z(n9566) );
  CAN2XL U16876 ( .A(n18017), .B(poly0_shifted[164]), .Z(n16995) );
  CANR1XL U16877 ( .A(Poly0[164]), .B(n17314), .C(n16995), .Z(n16996) );
  COND1XL U16878 ( .A(n17316), .B(n12005), .C(n16996), .Z(n9413) );
  CANR2X1 U16879 ( .A(n17750), .B(Poly8[73]), .C(n17266), .D(poly8_shifted[73]), .Z(n16997) );
  COND1XL U16880 ( .A(n12002), .B(n17750), .C(n16997), .Z(n11328) );
  CANR2X1 U16881 ( .A(n16694), .B(poly14_shifted[248]), .C(n17560), .D(
        poly14_shifted[232]), .Z(n16998) );
  COND1XL U16882 ( .A(n17166), .B(n16694), .C(n16998), .Z(n10173) );
  CANR2X1 U16883 ( .A(n16694), .B(poly14_shifted[262]), .C(n16999), .D(
        poly14_shifted[246]), .Z(n17000) );
  COND1XL U16884 ( .A(n17001), .B(n16694), .C(n17000), .Z(n10159) );
  CANR2X1 U16885 ( .A(n17969), .B(poly13_shifted[93]), .C(n17668), .D(
        poly13_shifted[79]), .Z(n17002) );
  COND1XL U16886 ( .A(n17196), .B(n17969), .C(n17002), .Z(n10981) );
  CANR2X1 U16887 ( .A(n17053), .B(poly1_shifted[233]), .C(n17965), .D(
        poly1_shifted[222]), .Z(n17003) );
  COND1XL U16888 ( .A(n17004), .B(n17053), .C(n17003), .Z(n9135) );
  CANR2XL U16889 ( .A(n12997), .B(poly12_shifted[26]), .C(n17215), .D(
        Poly12[121]), .Z(n17005) );
  COND1XL U16890 ( .A(n12014), .B(n12997), .C(n17005), .Z(n10522) );
  CANR2X1 U16891 ( .A(n17273), .B(poly7_shifted[219]), .C(n17552), .D(
        poly7_shifted[207]), .Z(n17006) );
  COND1XL U16892 ( .A(n17196), .B(n17273), .C(n17006), .Z(n9897) );
  CANR2X1 U16893 ( .A(n17987), .B(poly13_shifted[457]), .C(n17401), .D(
        poly13_shifted[443]), .Z(n17007) );
  COND1XL U16894 ( .A(n17741), .B(n17987), .C(n17007), .Z(n10617) );
  CANR2X1 U16895 ( .A(n13129), .B(Poly14[176]), .C(n16702), .D(
        poly14_shifted[176]), .Z(n17008) );
  COND1XL U16896 ( .A(n17211), .B(n13129), .C(n17008), .Z(n10229) );
  CANR2XL U16897 ( .A(n12958), .B(poly14_shifted[93]), .C(n17238), .D(
        poly14_shifted[77]), .Z(n17009) );
  COND1XL U16898 ( .A(n17090), .B(n12958), .C(n17009), .Z(n10328) );
  CANR2X1 U16899 ( .A(n17603), .B(poly13_shifted[351]), .C(n16919), .D(
        poly13_shifted[337]), .Z(n17010) );
  COND1XL U16900 ( .A(n17173), .B(n17603), .C(n17010), .Z(n10723) );
  CANR2XL U16901 ( .A(n13129), .B(poly14_shifted[179]), .C(n17285), .D(
        poly14_shifted[163]), .Z(n17011) );
  COND1XL U16902 ( .A(n13275), .B(n13129), .C(n17011), .Z(n10242) );
  CANR2X1 U16903 ( .A(n18002), .B(poly14_shifted[45]), .C(n17362), .D(
        poly14_shifted[29]), .Z(n17012) );
  COND1XL U16904 ( .A(n17185), .B(n18002), .C(n17012), .Z(n10376) );
  CANR2X1 U16905 ( .A(n12161), .B(Poly12[65]), .C(n17642), .D(
        poly12_shifted[65]), .Z(n17013) );
  COND1XL U16906 ( .A(n16950), .B(n12161), .C(n17013), .Z(n10467) );
  CANR2X1 U16907 ( .A(n17977), .B(Poly13[155]), .C(n17466), .D(
        poly13_shifted[155]), .Z(n17014) );
  COND1XL U16908 ( .A(n17741), .B(n17977), .C(n17014), .Z(n10905) );
  CANR2X1 U16909 ( .A(n17053), .B(poly1_shifted[231]), .C(n17504), .D(
        poly1_shifted[220]), .Z(n17015) );
  COND1XL U16910 ( .A(n11978), .B(n17053), .C(n17015), .Z(n9137) );
  CANR2XL U16911 ( .A(n12932), .B(poly14_shifted[286]), .C(n17136), .D(
        poly14_shifted[270]), .Z(n17017) );
  COND1XL U16912 ( .A(n12764), .B(n12932), .C(n17017), .Z(n10135) );
  CANR2X1 U16913 ( .A(n12008), .B(poly14_shifted[161]), .C(n17655), .D(
        poly14_shifted[145]), .Z(n17018) );
  COND1XL U16914 ( .A(n17173), .B(n12008), .C(n17018), .Z(n10260) );
  CANR2X1 U16915 ( .A(n17955), .B(poly9_shifted[77]), .C(n16488), .D(
        poly9_shifted[66]), .Z(n17019) );
  COND1XL U16916 ( .A(n16303), .B(n17955), .C(n17019), .Z(n11239) );
  CANR2X1 U16917 ( .A(n17332), .B(poly1_shifted[340]), .C(n16427), .D(
        poly1_shifted[329]), .Z(n17020) );
  COND1XL U16918 ( .A(n17208), .B(n17332), .C(n17020), .Z(n9028) );
  CANR2X1 U16919 ( .A(n17430), .B(Poly13[518]), .C(n17655), .D(
        poly13_shifted[518]), .Z(n17021) );
  COND1XL U16920 ( .A(n16779), .B(n17430), .C(n17021), .Z(n10542) );
  CANR2X1 U16921 ( .A(n17955), .B(poly9_shifted[81]), .C(n17105), .D(
        poly9_shifted[70]), .Z(n17022) );
  COND1XL U16922 ( .A(n17757), .B(n17955), .C(n17022), .Z(n11235) );
  CANR2X1 U16923 ( .A(n17990), .B(poly13_shifted[477]), .C(n17203), .D(
        poly13_shifted[463]), .Z(n17023) );
  COND1XL U16924 ( .A(n17196), .B(n17990), .C(n17023), .Z(n10597) );
  CANR2X1 U16925 ( .A(n17955), .B(poly9_shifted[75]), .C(n16985), .D(
        poly9_shifted[64]), .Z(n17024) );
  COND1XL U16926 ( .A(n12011), .B(n17955), .C(n17024), .Z(n11241) );
  CIVXL U16927 ( .A(n17675), .Z(n17025) );
  CANR2X1 U16928 ( .A(n12185), .B(poly11_shifted[18]), .C(n17209), .D(n17025), 
        .Z(n17026) );
  COND1XL U16929 ( .A(n13275), .B(n12185), .C(n17026), .Z(n11186) );
  CANR2XL U16930 ( .A(n18191), .B(poly1_shifted[283]), .C(n17998), .D(
        poly1_shifted[272]), .Z(n17027) );
  COND1XL U16931 ( .A(n17211), .B(n18191), .C(n17027), .Z(n9085) );
  CANR2X1 U16932 ( .A(n17982), .B(poly13_shifted[387]), .C(n16307), .D(
        poly13_shifted[373]), .Z(n17028) );
  COND1XL U16933 ( .A(n12006), .B(n17982), .C(n17028), .Z(n10687) );
  CANR2X1 U16934 ( .A(n18198), .B(poly1_shifted[299]), .C(n18047), .D(
        poly1_shifted[288]), .Z(n17029) );
  COND1XL U16935 ( .A(n12011), .B(n18198), .C(n17029), .Z(n9069) );
  CANR2X1 U16936 ( .A(n17595), .B(poly13_shifted[252]), .C(n17121), .D(
        poly13_shifted[238]), .Z(n17030) );
  COND1XL U16937 ( .A(n12764), .B(n17595), .C(n17030), .Z(n10822) );
  CANR2X1 U16938 ( .A(n12009), .B(poly14_shifted[122]), .C(n17449), .D(
        poly14_shifted[106]), .Z(n17032) );
  COND1XL U16939 ( .A(n12014), .B(n12009), .C(n17032), .Z(n10299) );
  CANR2X1 U16940 ( .A(n17491), .B(poly13_shifted[518]), .C(n17545), .D(
        poly13_shifted[504]), .Z(n17033) );
  COND1XL U16941 ( .A(n16179), .B(n17491), .C(n17033), .Z(n10556) );
  CANR2XL U16942 ( .A(n17430), .B(Poly13[515]), .C(n17206), .D(
        poly13_shifted[515]), .Z(n17034) );
  COND1XL U16943 ( .A(n13275), .B(n17430), .C(n17034), .Z(n10545) );
  CANR2X1 U16944 ( .A(n17731), .B(Poly9[21]), .C(n17655), .D(poly9_shifted[21]), .Z(n17035) );
  COND1XL U16945 ( .A(n17036), .B(n17731), .C(n17035), .Z(n11284) );
  CANR2X1 U16946 ( .A(n17500), .B(poly0_shifted[64]), .C(n17508), .D(
        poly0_shifted[46]), .Z(n17037) );
  COND1XL U16947 ( .A(n17502), .B(n17699), .C(n17037), .Z(n9531) );
  CANR2X1 U16948 ( .A(n17491), .B(poly13_shifted[511]), .C(n17533), .D(
        poly13_shifted[497]), .Z(n17038) );
  COND1XL U16949 ( .A(n17173), .B(n17491), .C(n17038), .Z(n10563) );
  CANR2X1 U16950 ( .A(n12012), .B(poly1_shifted[97]), .C(n16435), .D(
        poly1_shifted[86]), .Z(n17039) );
  COND1XL U16951 ( .A(n17753), .B(n12012), .C(n17039), .Z(n9271) );
  CANR2X1 U16952 ( .A(n12210), .B(poly1_shifted[196]), .C(n17398), .D(
        poly1_shifted[185]), .Z(n17040) );
  COND1XL U16953 ( .A(n17123), .B(n12210), .C(n17040), .Z(n9172) );
  CEOXL U16954 ( .A(Poly13[517]), .B(Poly13[390]), .Z(n17041) );
  CANR2X1 U16955 ( .A(n17043), .B(poly13_shifted[418]), .C(n17453), .D(n17041), 
        .Z(n17042) );
  COND1XL U16956 ( .A(n16391), .B(n17043), .C(n17042), .Z(n10656) );
  CANR2X1 U16957 ( .A(n17610), .B(poly1_shifted[139]), .C(n17099), .D(
        poly1_shifted[128]), .Z(n17044) );
  COND1XL U16958 ( .A(n12011), .B(n17610), .C(n17044), .Z(n9229) );
  CANR2X1 U16959 ( .A(n12012), .B(poly1_shifted[104]), .C(n17598), .D(
        poly1_shifted[93]), .Z(n17046) );
  COND1XL U16960 ( .A(n17185), .B(n12012), .C(n17046), .Z(n9264) );
  CIVXL U16961 ( .A(poly5_shifted[58]), .Z(n17049) );
  CANR2X1 U16962 ( .A(n17047), .B(n13028), .C(n16644), .D(poly5_shifted[44]), 
        .Z(n17048) );
  COND1XL U16963 ( .A(n17050), .B(n17049), .C(n17048), .Z(n11482) );
  CANR2X1 U16964 ( .A(n17603), .B(poly13_shifted[354]), .C(n16787), .D(
        poly13_shifted[340]), .Z(n17051) );
  COND1XL U16965 ( .A(n16391), .B(n17603), .C(n17051), .Z(n10720) );
  CANR2X1 U16966 ( .A(n17053), .B(poly1_shifted[203]), .C(n16372), .D(
        poly1_shifted[192]), .Z(n17052) );
  COND1XL U16967 ( .A(n12011), .B(n17053), .C(n17052), .Z(n9165) );
  CANR2X1 U16968 ( .A(n16425), .B(poly1_shifted[114]), .C(n16479), .D(
        poly1_shifted[103]), .Z(n17054) );
  COND1XL U16969 ( .A(n16939), .B(n16425), .C(n17054), .Z(n9254) );
  CANR2X1 U16970 ( .A(n17990), .B(poly13_shifted[471]), .C(n16540), .D(
        poly13_shifted[457]), .Z(n17055) );
  COND1XL U16971 ( .A(n12002), .B(n17990), .C(n17055), .Z(n10603) );
  CANR2X1 U16972 ( .A(n17503), .B(Poly0[10]), .C(n17198), .D(Poly0[212]), .Z(
        n17056) );
  COND1XL U16973 ( .A(n17506), .B(n12014), .C(n17056), .Z(n9567) );
  CANR2X1 U16974 ( .A(n17671), .B(Poly0[150]), .C(n17527), .D(
        poly0_shifted[150]), .Z(n17057) );
  COND1XL U16975 ( .A(n17674), .B(n17753), .C(n17057), .Z(n9427) );
  CANR2X1 U16976 ( .A(n17969), .B(poly13_shifted[81]), .C(n17178), .D(
        poly13_shifted[67]), .Z(n17058) );
  COND1XL U16977 ( .A(n13275), .B(n17969), .C(n17058), .Z(n10993) );
  CANR2X1 U16978 ( .A(n17595), .B(poly13_shifted[265]), .C(n17280), .D(
        poly13_shifted[251]), .Z(n17059) );
  COND1XL U16979 ( .A(n17741), .B(n17595), .C(n17059), .Z(n10809) );
  CANR2XL U16980 ( .A(n16695), .B(poly0_shifted[22]), .C(n17503), .D(Poly0[22]), .Z(n17060) );
  COND1XL U16981 ( .A(n17506), .B(n17753), .C(n17060), .Z(n9555) );
  CANR2XL U16982 ( .A(n17552), .B(Poly0[218]), .C(n17503), .D(Poly0[16]), .Z(
        n17061) );
  COND1XL U16983 ( .A(n17506), .B(n17062), .C(n17061), .Z(n9561) );
  CANR2X1 U16984 ( .A(n17063), .B(Poly0[215]), .C(n17503), .D(Poly0[13]), .Z(
        n17064) );
  COND1XL U16985 ( .A(n17506), .B(n17065), .C(n17064), .Z(n9564) );
  CANR2X1 U16986 ( .A(n17209), .B(Poly0[217]), .C(n17503), .D(Poly0[15]), .Z(
        n17066) );
  COND1XL U16987 ( .A(n17506), .B(n17196), .C(n17066), .Z(n9562) );
  CANR2X1 U16988 ( .A(n17466), .B(Poly0[211]), .C(n17503), .D(Poly0[9]), .Z(
        n17067) );
  COND1XL U16989 ( .A(n17506), .B(n17208), .C(n17067), .Z(n9568) );
  CANR2XL U16990 ( .A(n17280), .B(Poly0[206]), .C(n17503), .D(
        poly0_shifted[22]), .Z(n17068) );
  COND1XL U16991 ( .A(n17506), .B(n12005), .C(n17068), .Z(n9573) );
  CANR2XL U16992 ( .A(n17063), .B(Poly0[203]), .C(n17503), .D(
        poly0_shifted[19]), .Z(n17069) );
  COND1XL U16993 ( .A(n17506), .B(n17711), .C(n17069), .Z(n9576) );
  CANR2X1 U16994 ( .A(n16307), .B(Poly0[216]), .C(n17503), .D(Poly0[14]), .Z(
        n17070) );
  COND1XL U16995 ( .A(n17506), .B(n17699), .C(n17070), .Z(n9563) );
  CANR2XL U16996 ( .A(n17288), .B(Poly0[205]), .C(n17503), .D(
        poly0_shifted[21]), .Z(n17071) );
  COND1XL U16997 ( .A(n17506), .B(n13275), .C(n17071), .Z(n9574) );
  CANR2X1 U16998 ( .A(n17072), .B(Poly0[214]), .C(n17503), .D(Poly0[12]), .Z(
        n17073) );
  COND1XL U16999 ( .A(n17506), .B(n17087), .C(n17073), .Z(n9565) );
  CANR2XL U17000 ( .A(n17280), .B(Poly0[209]), .C(n17503), .D(Poly0[7]), .Z(
        n17074) );
  COND1XL U17001 ( .A(n17506), .B(n17718), .C(n17074), .Z(n9570) );
  CANR2X1 U17002 ( .A(n17965), .B(Poly0[219]), .C(n17503), .D(Poly0[17]), .Z(
        n17075) );
  COND1XL U17003 ( .A(n17506), .B(n17076), .C(n17075), .Z(n9560) );
  CANR2X1 U17004 ( .A(n17533), .B(poly0_shifted[59]), .C(n17500), .D(
        poly0_shifted[77]), .Z(n17077) );
  COND1XL U17005 ( .A(n17502), .B(n17741), .C(n17077), .Z(n9518) );
  CANR2X1 U17006 ( .A(n16435), .B(poly0_shifted[190]), .C(poly0_shifted[208]), 
        .D(n17314), .Z(n17078) );
  COND1XL U17007 ( .A(n17316), .B(n17004), .C(n17078), .Z(n9387) );
  CANR2X1 U17008 ( .A(n17398), .B(poly0_shifted[149]), .C(n17671), .D(
        poly0_shifted[167]), .Z(n17079) );
  COND1XL U17009 ( .A(n17674), .B(n12006), .C(n17079), .Z(n9428) );
  CANR2X1 U17010 ( .A(n12401), .B(Poly7[400]), .C(n17488), .D(
        poly7_shifted[400]), .Z(n17080) );
  COND1XL U17011 ( .A(n17211), .B(n12401), .C(n17080), .Z(n9704) );
  CANR2X1 U17012 ( .A(n12401), .B(poly7_shifted[407]), .C(n17105), .D(
        poly7_shifted[395]), .Z(n17081) );
  COND1XL U17013 ( .A(n16994), .B(n12401), .C(n17081), .Z(n9709) );
  CANR2X1 U17014 ( .A(n12401), .B(Poly7[409]), .C(n17099), .D(
        poly7_shifted[409]), .Z(n17082) );
  COND1XL U17015 ( .A(n17123), .B(n12401), .C(n17082), .Z(n9695) );
  CANR2X1 U17016 ( .A(n12401), .B(poly7_shifted[397]), .C(n17535), .D(
        poly7_shifted[385]), .Z(n17083) );
  COND1XL U17017 ( .A(n17697), .B(n12401), .C(n17083), .Z(n9719) );
  CANR2X1 U17018 ( .A(n12401), .B(poly7_shifted[405]), .C(n17121), .D(
        poly7_shifted[393]), .Z(n17084) );
  COND1XL U17019 ( .A(n17208), .B(n12401), .C(n17084), .Z(n9711) );
  CANR2XL U17020 ( .A(n12401), .B(Poly7[408]), .C(n17535), .D(
        poly7_shifted[408]), .Z(n17085) );
  COND1XL U17021 ( .A(n16179), .B(n12401), .C(n17085), .Z(n9696) );
  CANR2X1 U17022 ( .A(n12401), .B(poly7_shifted[408]), .C(n17535), .D(
        poly7_shifted[396]), .Z(n17086) );
  COND1XL U17023 ( .A(n17087), .B(n12401), .C(n17086), .Z(n9708) );
  CANR2X1 U17024 ( .A(n12401), .B(Poly7[399]), .C(n17634), .D(
        poly7_shifted[399]), .Z(n17088) );
  COND1XL U17025 ( .A(n17196), .B(n12401), .C(n17088), .Z(n9705) );
  CANR2X1 U17026 ( .A(n12401), .B(poly7_shifted[409]), .C(n17535), .D(
        poly7_shifted[397]), .Z(n17089) );
  COND1XL U17027 ( .A(n17090), .B(n12401), .C(n17089), .Z(n9707) );
  CANR2X1 U17028 ( .A(n12401), .B(poly7_shifted[396]), .C(n17535), .D(
        poly7_shifted[384]), .Z(n17091) );
  COND1XL U17029 ( .A(n12011), .B(n12401), .C(n17091), .Z(n9720) );
  CANR2X1 U17030 ( .A(n12401), .B(poly7_shifted[404]), .C(n17390), .D(
        poly7_shifted[392]), .Z(n17092) );
  COND1XL U17031 ( .A(n17166), .B(n12401), .C(n17092), .Z(n9712) );
  CANR2X1 U17032 ( .A(n12401), .B(poly7_shifted[399]), .C(n17453), .D(
        poly7_shifted[387]), .Z(n17093) );
  COND1XL U17033 ( .A(n13275), .B(n12401), .C(n17093), .Z(n9717) );
  CANR2X1 U17034 ( .A(n17094), .B(Poly0[202]), .C(n17503), .D(
        poly0_shifted[18]), .Z(n17095) );
  COND1XL U17035 ( .A(n17506), .B(n17751), .C(n17095), .Z(n9577) );
  CANR2XL U17036 ( .A(n18234), .B(poly0_shifted[21]), .C(n17503), .D(Poly0[21]), .Z(n17096) );
  COND1XL U17037 ( .A(n17506), .B(n12006), .C(n17096), .Z(n9556) );
  CANR2X1 U17038 ( .A(n12170), .B(poly7_shifted[57]), .C(n17453), .D(
        poly7_shifted[45]), .Z(n17097) );
  COND1XL U17039 ( .A(n17065), .B(n12170), .C(n17097), .Z(n10059) );
  CANR2X1 U17040 ( .A(n12170), .B(poly7_shifted[58]), .C(n17552), .D(
        poly7_shifted[46]), .Z(n17098) );
  COND1XL U17041 ( .A(n17699), .B(n12170), .C(n17098), .Z(n10058) );
  CANR2X1 U17042 ( .A(n12170), .B(Poly7[53]), .C(n17099), .D(poly7_shifted[53]), .Z(n17100) );
  COND1XL U17043 ( .A(n12006), .B(n12170), .C(n17100), .Z(n10051) );
  CANR2X1 U17044 ( .A(n12170), .B(Poly7[57]), .C(n17206), .D(poly7_shifted[57]), .Z(n17101) );
  COND1XL U17045 ( .A(n17123), .B(n12170), .C(n17101), .Z(n10047) );
  CANR2X1 U17046 ( .A(n12170), .B(poly7_shifted[56]), .C(n17965), .D(
        poly7_shifted[44]), .Z(n17102) );
  COND1XL U17047 ( .A(n17087), .B(n12170), .C(n17102), .Z(n10060) );
  CANR2X1 U17048 ( .A(n12170), .B(Poly7[59]), .C(n17398), .D(poly7_shifted[59]), .Z(n17103) );
  COND1XL U17049 ( .A(n17741), .B(n12170), .C(n17103), .Z(n10045) );
  CANR2X1 U17050 ( .A(n12170), .B(Poly7[56]), .C(n17203), .D(poly7_shifted[56]), .Z(n17104) );
  COND1XL U17051 ( .A(n17721), .B(n12170), .C(n17104), .Z(n10048) );
  CANR2X1 U17052 ( .A(n12170), .B(Poly7[48]), .C(n17105), .D(poly7_shifted[48]), .Z(n17106) );
  COND1XL U17053 ( .A(n17211), .B(n12170), .C(n17106), .Z(n10056) );
  CANR2X1 U17054 ( .A(n12170), .B(poly7_shifted[55]), .C(n16787), .D(
        poly7_shifted[43]), .Z(n17107) );
  COND1XL U17055 ( .A(n16994), .B(n12170), .C(n17107), .Z(n10061) );
  CANR2X1 U17056 ( .A(n12170), .B(Poly7[54]), .C(n17198), .D(poly7_shifted[54]), .Z(n17108) );
  COND1XL U17057 ( .A(n17753), .B(n12170), .C(n17108), .Z(n10050) );
  CANR2X1 U17058 ( .A(n12170), .B(Poly7[49]), .C(n16435), .D(poly7_shifted[49]), .Z(n17109) );
  COND1XL U17059 ( .A(n17173), .B(n12170), .C(n17109), .Z(n10055) );
  CEOXL U17060 ( .A(Poly7[400]), .B(Poly7[49]), .Z(n17110) );
  CANR2X1 U17061 ( .A(n12170), .B(poly7_shifted[73]), .C(n17198), .D(n17110), 
        .Z(n17111) );
  COND1XL U17062 ( .A(n17185), .B(n12170), .C(n17111), .Z(n10043) );
  CANR2X1 U17063 ( .A(n12170), .B(poly7_shifted[59]), .C(n16695), .D(
        poly7_shifted[47]), .Z(n17112) );
  COND1XL U17064 ( .A(n17196), .B(n12170), .C(n17112), .Z(n10057) );
  CANR2X1 U17065 ( .A(n13040), .B(poly7_shifted[333]), .C(n17449), .D(
        poly7_shifted[321]), .Z(n17113) );
  COND1XL U17066 ( .A(n17697), .B(n13040), .C(n17113), .Z(n9783) );
  CANR2X1 U17067 ( .A(n13040), .B(poly7_shifted[335]), .C(n17545), .D(
        poly7_shifted[323]), .Z(n17114) );
  COND1XL U17068 ( .A(n13275), .B(n13040), .C(n17114), .Z(n9781) );
  CANR2X1 U17069 ( .A(n13040), .B(poly7_shifted[332]), .C(n17105), .D(
        poly7_shifted[320]), .Z(n17115) );
  COND1XL U17070 ( .A(n12011), .B(n13040), .C(n17115), .Z(n9784) );
  CANR2X1 U17071 ( .A(n13040), .B(poly7_shifted[340]), .C(n17552), .D(
        poly7_shifted[328]), .Z(n17116) );
  COND1XL U17072 ( .A(n17166), .B(n13040), .C(n17116), .Z(n9776) );
  CANR2X1 U17073 ( .A(n13040), .B(poly7_shifted[353]), .C(n17136), .D(
        poly7_shifted[341]), .Z(n17117) );
  COND1XL U17074 ( .A(n12006), .B(n13040), .C(n17117), .Z(n9763) );
  CANR2X1 U17075 ( .A(n13040), .B(poly7_shifted[338]), .C(n17642), .D(
        poly7_shifted[326]), .Z(n17118) );
  COND1XL U17076 ( .A(n16779), .B(n13040), .C(n17118), .Z(n9778) );
  CANR2X1 U17077 ( .A(n13040), .B(poly7_shifted[345]), .C(n17401), .D(
        poly7_shifted[333]), .Z(n17119) );
  COND1XL U17078 ( .A(n17090), .B(n13040), .C(n17119), .Z(n9771) );
  CANR2X1 U17079 ( .A(n13040), .B(poly7_shifted[362]), .C(n17504), .D(
        poly7_shifted[350]), .Z(n17120) );
  COND1XL U17080 ( .A(n17004), .B(n13040), .C(n17120), .Z(n9754) );
  CANR2X1 U17081 ( .A(n13040), .B(poly7_shifted[357]), .C(n17121), .D(
        poly7_shifted[345]), .Z(n17122) );
  COND1XL U17082 ( .A(n17123), .B(n13040), .C(n17122), .Z(n9759) );
  CEOXL U17083 ( .A(Poly3[72]), .B(Poly3[80]), .Z(n17124) );
  CENX1 U17084 ( .A(Poly3[47]), .B(n17124), .Z(n17125) );
  CNR2XL U17085 ( .A(n17826), .B(n17125), .Z(n17126) );
  CANR1XL U17086 ( .A(poly3_shifted[75]), .B(n17587), .C(n17126), .Z(n17127)
         );
  COND1XL U17087 ( .A(n17185), .B(n17589), .C(n17127), .Z(n8879) );
  CANR2X1 U17088 ( .A(n18028), .B(poly7_shifted[322]), .C(n17295), .D(
        poly7_shifted[310]), .Z(n17128) );
  COND1XL U17089 ( .A(n17753), .B(n18028), .C(n17128), .Z(n9794) );
  CANR2X1 U17090 ( .A(n18028), .B(poly7_shifted[331]), .C(n17598), .D(
        poly7_shifted[319]), .Z(n17129) );
  COND1XL U17091 ( .A(n17188), .B(n18028), .C(n17129), .Z(n9785) );
  CANR2X1 U17092 ( .A(n18028), .B(poly7_shifted[321]), .C(n16502), .D(
        poly7_shifted[309]), .Z(n17130) );
  COND1XL U17093 ( .A(n12006), .B(n18028), .C(n17130), .Z(n9795) );
  CANR2X1 U17094 ( .A(n18028), .B(poly7_shifted[316]), .C(n17449), .D(
        poly7_shifted[304]), .Z(n17131) );
  COND1XL U17095 ( .A(n17211), .B(n18028), .C(n17131), .Z(n9800) );
  CANR2X1 U17096 ( .A(n18028), .B(poly7_shifted[328]), .C(n17545), .D(
        poly7_shifted[316]), .Z(n17132) );
  COND1XL U17097 ( .A(n11978), .B(n18028), .C(n17132), .Z(n9788) );
  CANR2X1 U17098 ( .A(n18028), .B(poly7_shifted[305]), .C(n17136), .D(
        poly7_shifted[293]), .Z(n17133) );
  COND1XL U17099 ( .A(n11985), .B(n18028), .C(n17133), .Z(n9811) );
  CANR2X1 U17100 ( .A(n18028), .B(poly7_shifted[312]), .C(n17535), .D(
        poly7_shifted[300]), .Z(n17134) );
  COND1XL U17101 ( .A(n17218), .B(n18028), .C(n17134), .Z(n9804) );
  CANR2X1 U17102 ( .A(n18028), .B(poly7_shifted[308]), .C(n16323), .D(
        poly7_shifted[296]), .Z(n17135) );
  COND1XL U17103 ( .A(n17166), .B(n18028), .C(n17135), .Z(n9808) );
  CANR2X1 U17104 ( .A(n13040), .B(poly7_shifted[341]), .C(n17136), .D(
        poly7_shifted[329]), .Z(n17137) );
  COND1XL U17105 ( .A(n17208), .B(n13040), .C(n17137), .Z(n9775) );
  CANR2X1 U17106 ( .A(n13040), .B(poly7_shifted[344]), .C(n17203), .D(
        poly7_shifted[332]), .Z(n17138) );
  COND1XL U17107 ( .A(n17087), .B(n13040), .C(n17138), .Z(n9772) );
  CANR2X1 U17108 ( .A(n13040), .B(poly7_shifted[346]), .C(n17295), .D(
        poly7_shifted[334]), .Z(n17139) );
  COND1XL U17109 ( .A(n12764), .B(n13040), .C(n17139), .Z(n9770) );
  CANR2X1 U17110 ( .A(n13040), .B(poly7_shifted[356]), .C(n16985), .D(
        poly7_shifted[344]), .Z(n17140) );
  COND1XL U17111 ( .A(n16179), .B(n13040), .C(n17140), .Z(n9760) );
  CANR2X1 U17112 ( .A(n13040), .B(poly7_shifted[354]), .C(n17545), .D(
        poly7_shifted[342]), .Z(n17141) );
  COND1XL U17113 ( .A(n17753), .B(n13040), .C(n17141), .Z(n9762) );
  CANR2X1 U17114 ( .A(n13040), .B(poly7_shifted[334]), .C(n17295), .D(
        poly7_shifted[322]), .Z(n17142) );
  COND1XL U17115 ( .A(n16775), .B(n13040), .C(n17142), .Z(n9782) );
  CANR2X1 U17116 ( .A(n17587), .B(Poly3[40]), .C(n17245), .D(poly3_shifted[40]), .Z(n17143) );
  COND1XL U17117 ( .A(n17163), .B(n17589), .C(n17143), .Z(n8900) );
  CANR2X1 U17118 ( .A(n17587), .B(Poly3[32]), .C(n17144), .D(poly3_shifted[32]), .Z(n17145) );
  COND1XL U17119 ( .A(n17751), .B(n17262), .C(n17145), .Z(n8908) );
  CANR2X1 U17120 ( .A(n17587), .B(Poly3[39]), .C(n16540), .D(poly3_shifted[39]), .Z(n17146) );
  COND1XL U17121 ( .A(n16939), .B(n17589), .C(n17146), .Z(n8901) );
  CANR2X1 U17122 ( .A(n17587), .B(Poly3[44]), .C(n17356), .D(poly3_shifted[44]), .Z(n17147) );
  COND1XL U17123 ( .A(n17087), .B(n17589), .C(n17147), .Z(n8896) );
  CANR2X1 U17124 ( .A(n17587), .B(Poly3[35]), .C(n17266), .D(poly3_shifted[35]), .Z(n17148) );
  COND1XL U17125 ( .A(n13275), .B(n17589), .C(n17148), .Z(n8905) );
  CANR2X1 U17126 ( .A(n17587), .B(Poly3[43]), .C(n17245), .D(poly3_shifted[43]), .Z(n17149) );
  COND1XL U17127 ( .A(n16994), .B(n17589), .C(n17149), .Z(n8897) );
  CENX1 U17128 ( .A(Poly3[70]), .B(Poly3[78]), .Z(n17150) );
  CENX1 U17129 ( .A(Poly3[45]), .B(n17150), .Z(n17151) );
  CANR2X1 U17130 ( .A(n17587), .B(poly3_shifted[73]), .C(n17158), .D(n17151), 
        .Z(n17152) );
  COND1XL U17131 ( .A(n17741), .B(n17587), .C(n17152), .Z(n8881) );
  CANR2X1 U17132 ( .A(n17587), .B(Poly3[33]), .C(n17523), .D(poly3_shifted[33]), .Z(n17153) );
  COND1XL U17133 ( .A(n17697), .B(n17589), .C(n17153), .Z(n8907) );
  CANR2X1 U17134 ( .A(n17587), .B(Poly3[37]), .C(n17245), .D(poly3_shifted[37]), .Z(n17154) );
  COND1XL U17135 ( .A(n11987), .B(n17589), .C(n17154), .Z(n8903) );
  CANR2X1 U17136 ( .A(n17587), .B(Poly3[38]), .C(n17156), .D(poly3_shifted[38]), .Z(n17155) );
  COND1XL U17137 ( .A(n16779), .B(n17589), .C(n17155), .Z(n8902) );
  CANR2X1 U17138 ( .A(n17587), .B(Poly3[41]), .C(n17156), .D(poly3_shifted[41]), .Z(n17157) );
  COND1XL U17139 ( .A(n17208), .B(n17589), .C(n17157), .Z(n8899) );
  CANR2X1 U17140 ( .A(n17587), .B(Poly3[34]), .C(n17158), .D(poly3_shifted[34]), .Z(n17159) );
  COND1XL U17141 ( .A(n16775), .B(n17262), .C(n17159), .Z(n8906) );
  CNR2IXL U17142 ( .B(poly7_shifted[104]), .A(n17160), .Z(n17161) );
  CANR1XL U17143 ( .A(poly7_shifted[116]), .B(n17217), .C(n17161), .Z(n17162)
         );
  COND1XL U17144 ( .A(n17163), .B(n17217), .C(n17162), .Z(n10000) );
  CANR2X1 U17145 ( .A(n13070), .B(poly7_shifted[146]), .C(n17290), .D(
        poly7_shifted[134]), .Z(n17164) );
  COND1XL U17146 ( .A(n17757), .B(n13070), .C(n17164), .Z(n9970) );
  CANR2X1 U17147 ( .A(n13070), .B(poly7_shifted[148]), .C(n17209), .D(
        poly7_shifted[136]), .Z(n17165) );
  COND1XL U17148 ( .A(n17166), .B(n13070), .C(n17165), .Z(n9968) );
  CANR2X1 U17149 ( .A(n13070), .B(poly7_shifted[157]), .C(n17178), .D(
        poly7_shifted[145]), .Z(n17167) );
  COND1XL U17150 ( .A(n17173), .B(n13070), .C(n17167), .Z(n9959) );
  CANR2X1 U17151 ( .A(n12401), .B(\dataselector_shifted[0] ), .C(n17390), .D(
        poly7_shifted[404]), .Z(n17168) );
  COND1XL U17152 ( .A(n16391), .B(n12401), .C(n17168), .Z(n9700) );
  CANR2X1 U17153 ( .A(n12401), .B(Poly7[406]), .C(n17203), .D(
        poly7_shifted[406]), .Z(n17169) );
  COND1XL U17154 ( .A(n17753), .B(n12401), .C(n17169), .Z(n9698) );
  CANR2X1 U17155 ( .A(n12401), .B(poly7_shifted[406]), .C(n16985), .D(
        poly7_shifted[394]), .Z(n17170) );
  COND1XL U17156 ( .A(n12014), .B(n12401), .C(n17170), .Z(n9710) );
  CANR2X1 U17157 ( .A(n12401), .B(Poly7[405]), .C(n17398), .D(
        poly7_shifted[405]), .Z(n17171) );
  COND1XL U17158 ( .A(n12006), .B(n12401), .C(n17171), .Z(n9699) );
  CANR2X1 U17159 ( .A(n12401), .B(Poly7[401]), .C(n17174), .D(
        poly7_shifted[401]), .Z(n17172) );
  COND1XL U17160 ( .A(n17173), .B(n12401), .C(n17172), .Z(n9703) );
  CANR2X1 U17161 ( .A(n12401), .B(poly7_shifted[401]), .C(n17174), .D(
        poly7_shifted[389]), .Z(n17175) );
  COND1XL U17162 ( .A(n11983), .B(n12401), .C(n17175), .Z(n9715) );
  CANR2X1 U17163 ( .A(n12401), .B(poly7_shifted[410]), .C(n17998), .D(
        poly7_shifted[398]), .Z(n17176) );
  COND1XL U17164 ( .A(n12764), .B(n12401), .C(n17176), .Z(n9706) );
  CANR2X1 U17165 ( .A(n12401), .B(poly7_shifted[398]), .C(n17266), .D(
        poly7_shifted[386]), .Z(n17177) );
  COND1XL U17166 ( .A(n16303), .B(n12401), .C(n17177), .Z(n9718) );
  CANR2X1 U17167 ( .A(n13070), .B(poly7_shifted[145]), .C(n17178), .D(
        poly7_shifted[133]), .Z(n17179) );
  COND1XL U17168 ( .A(n11985), .B(n13070), .C(n17179), .Z(n9971) );
  CANR2X1 U17169 ( .A(n13070), .B(poly7_shifted[155]), .C(n17535), .D(
        poly7_shifted[143]), .Z(n17180) );
  COND1XL U17170 ( .A(n17196), .B(n13070), .C(n17180), .Z(n9961) );
  CANR2X1 U17171 ( .A(n13070), .B(poly7_shifted[150]), .C(n16787), .D(
        poly7_shifted[138]), .Z(n17181) );
  COND1XL U17172 ( .A(n12014), .B(n13070), .C(n17181), .Z(n9966) );
  CANR2X1 U17173 ( .A(n17217), .B(poly7_shifted[130]), .C(n17504), .D(
        poly7_shifted[118]), .Z(n17182) );
  COND1XL U17174 ( .A(n17753), .B(n17217), .C(n17182), .Z(n9986) );
  CANR2X1 U17175 ( .A(n17217), .B(poly7_shifted[118]), .C(n17965), .D(
        poly7_shifted[106]), .Z(n17183) );
  COND1XL U17176 ( .A(n12014), .B(n17217), .C(n17183), .Z(n9998) );
  CANR2X1 U17177 ( .A(n17217), .B(poly7_shifted[137]), .C(n17352), .D(
        poly7_shifted[125]), .Z(n17184) );
  COND1XL U17178 ( .A(n17185), .B(n17217), .C(n17184), .Z(n9979) );
  CANR2X1 U17179 ( .A(n17217), .B(poly7_shifted[125]), .C(n17352), .D(
        poly7_shifted[113]), .Z(n17186) );
  COND1XL U17180 ( .A(n17173), .B(n17217), .C(n17186), .Z(n9991) );
  CANR2X1 U17181 ( .A(n17217), .B(poly7_shifted[139]), .C(n17266), .D(
        poly7_shifted[127]), .Z(n17187) );
  COND1XL U17182 ( .A(n17188), .B(n17217), .C(n17187), .Z(n9977) );
  CANR2X1 U17183 ( .A(n17217), .B(poly7_shifted[111]), .C(n17063), .D(
        poly7_shifted[99]), .Z(n17189) );
  COND1XL U17184 ( .A(n13275), .B(n17217), .C(n17189), .Z(n10005) );
  CANR2X1 U17185 ( .A(n17217), .B(poly7_shifted[113]), .C(n17266), .D(
        poly7_shifted[101]), .Z(n17190) );
  COND1XL U17186 ( .A(n11987), .B(n17217), .C(n17190), .Z(n10003) );
  CANR2X1 U17187 ( .A(n17217), .B(poly7_shifted[109]), .C(n17198), .D(
        poly7_shifted[97]), .Z(n17191) );
  COND1XL U17188 ( .A(n16950), .B(n17217), .C(n17191), .Z(n10007) );
  CANR2X1 U17189 ( .A(n17217), .B(poly7_shifted[135]), .C(n16985), .D(
        poly7_shifted[123]), .Z(n17192) );
  COND1XL U17190 ( .A(n17741), .B(n17217), .C(n17192), .Z(n9981) );
  CANR2X1 U17191 ( .A(n17217), .B(poly7_shifted[121]), .C(n17198), .D(
        poly7_shifted[109]), .Z(n17193) );
  COND1XL U17192 ( .A(n17090), .B(n17217), .C(n17193), .Z(n9995) );
  CANR2X1 U17193 ( .A(n17217), .B(poly7_shifted[128]), .C(n16702), .D(
        poly7_shifted[116]), .Z(n17194) );
  COND1XL U17194 ( .A(n17707), .B(n17217), .C(n17194), .Z(n9988) );
  CANR2X1 U17195 ( .A(n17217), .B(poly7_shifted[123]), .C(n17458), .D(
        poly7_shifted[111]), .Z(n17195) );
  COND1XL U17196 ( .A(n17196), .B(n17217), .C(n17195), .Z(n9993) );
  CANR2X1 U17197 ( .A(n17217), .B(poly7_shifted[136]), .C(n17209), .D(
        poly7_shifted[124]), .Z(n17197) );
  COND1XL U17198 ( .A(n11978), .B(n17217), .C(n17197), .Z(n9980) );
  CANR2X1 U17199 ( .A(n17217), .B(poly7_shifted[133]), .C(n17198), .D(
        poly7_shifted[121]), .Z(n17199) );
  COND1XL U17200 ( .A(n17200), .B(n17217), .C(n17199), .Z(n9983) );
  CANR2X1 U17201 ( .A(n17217), .B(poly7_shifted[138]), .C(n17458), .D(
        poly7_shifted[126]), .Z(n17201) );
  COND1XL U17202 ( .A(n17004), .B(n17217), .C(n17201), .Z(n9978) );
  CANR2X1 U17203 ( .A(n17217), .B(poly7_shifted[110]), .C(n17203), .D(
        poly7_shifted[98]), .Z(n17202) );
  COND1XL U17204 ( .A(n16775), .B(n17217), .C(n17202), .Z(n10006) );
  CANR2X1 U17205 ( .A(n17217), .B(poly7_shifted[122]), .C(n17203), .D(
        poly7_shifted[110]), .Z(n17204) );
  COND1XL U17206 ( .A(n12764), .B(n17217), .C(n17204), .Z(n9994) );
  CANR2X1 U17207 ( .A(n17217), .B(poly7_shifted[129]), .C(n17206), .D(
        poly7_shifted[117]), .Z(n17205) );
  COND1XL U17208 ( .A(n12006), .B(n17217), .C(n17205), .Z(n9987) );
  CANR2X1 U17209 ( .A(n17217), .B(poly7_shifted[117]), .C(n17206), .D(
        poly7_shifted[105]), .Z(n17207) );
  COND1XL U17210 ( .A(n17208), .B(n17217), .C(n17207), .Z(n9999) );
  CANR2X1 U17211 ( .A(n17217), .B(poly7_shifted[124]), .C(n17209), .D(
        poly7_shifted[112]), .Z(n17210) );
  COND1XL U17212 ( .A(n17211), .B(n17217), .C(n17210), .Z(n9992) );
  CANR2X1 U17213 ( .A(n17217), .B(poly7_shifted[132]), .C(n17215), .D(
        poly7_shifted[120]), .Z(n17212) );
  COND1XL U17214 ( .A(n16179), .B(n17217), .C(n17212), .Z(n9984) );
  CANR2X1 U17215 ( .A(n17217), .B(poly7_shifted[108]), .C(n17215), .D(
        poly7_shifted[96]), .Z(n17213) );
  COND1XL U17216 ( .A(n12011), .B(n17217), .C(n17213), .Z(n10008) );
  CANR2X1 U17217 ( .A(n17217), .B(poly7_shifted[119]), .C(n17535), .D(
        poly7_shifted[107]), .Z(n17214) );
  COND1XL U17218 ( .A(n16994), .B(n17217), .C(n17214), .Z(n9997) );
  CANR2X1 U17219 ( .A(n17217), .B(poly7_shifted[120]), .C(n17215), .D(
        poly7_shifted[108]), .Z(n17216) );
  COND1XL U17220 ( .A(n17218), .B(n17217), .C(n17216), .Z(n9996) );
  CIVX1 U17221 ( .A(n17219), .Z(n17220) );
  CANR2X1 U17222 ( .A(n17220), .B(n17099), .C(poly4_shifted[20]), .D(n18230), 
        .Z(n17221) );
  COND1XL U17223 ( .A(n13275), .B(n18230), .C(n17221), .Z(n8853) );
  CEOXL U17224 ( .A(Poly4[43]), .B(Poly4[52]), .Z(n17223) );
  CENX1 U17225 ( .A(Poly4[51]), .B(Poly4[53]), .Z(n17222) );
  CENX1 U17226 ( .A(n17223), .B(n17222), .Z(n17224) );
  CENX1 U17227 ( .A(n17225), .B(n17224), .Z(n17226) );
  CENX1 U17228 ( .A(n17326), .B(n17226), .Z(n17227) );
  CNR2XL U17229 ( .A(n17227), .B(n17959), .Z(n17228) );
  CANR1XL U17230 ( .A(Poly4[60]), .B(n12153), .C(n17228), .Z(n17229) );
  COND1XL U17231 ( .A(n11978), .B(n12153), .C(n17229), .Z(n8796) );
  CANR2X1 U17232 ( .A(n17974), .B(poly13_shifted[115]), .C(n17755), .D(
        poly13_shifted[101]), .Z(n17230) );
  COND1XL U17233 ( .A(n11993), .B(n17974), .C(n17230), .Z(n10959) );
  CANR2X1 U17234 ( .A(n17430), .B(Poly13[517]), .C(n18047), .D(
        poly13_shifted[517]), .Z(n17231) );
  COND1XL U17235 ( .A(n11991), .B(n17430), .C(n17231), .Z(n10543) );
  CANR2X1 U17236 ( .A(n17491), .B(poly13_shifted[499]), .C(n16695), .D(
        poly13_shifted[485]), .Z(n17232) );
  COND1XL U17237 ( .A(n11981), .B(n17491), .C(n17232), .Z(n10575) );
  CEOXL U17238 ( .A(n17233), .B(Poly11[22]), .Z(n17234) );
  CANR2X1 U17239 ( .A(n17683), .B(Poly11[37]), .C(n17362), .D(n17234), .Z(
        n17235) );
  COND1XL U17240 ( .A(n11987), .B(n17747), .C(n17235), .Z(n11152) );
  CANR2X1 U17241 ( .A(n17667), .B(poly13_shifted[211]), .C(n17538), .D(
        poly13_shifted[197]), .Z(n17236) );
  COND1XL U17242 ( .A(n11983), .B(n17667), .C(n17236), .Z(n10863) );
  CANR2X1 U17243 ( .A(n17603), .B(poly13_shifted[339]), .C(n16326), .D(
        poly13_shifted[325]), .Z(n17237) );
  COND1XL U17244 ( .A(n11991), .B(n17603), .C(n17237), .Z(n10735) );
  CANR2X1 U17245 ( .A(n12206), .B(poly7_shifted[390]), .C(n17238), .D(
        poly7_shifted[378]), .Z(n17239) );
  COND1XL U17246 ( .A(n17735), .B(n12206), .C(n17239), .Z(n9726) );
  CANR2X1 U17247 ( .A(n17471), .B(poly7_shifted[102]), .C(n17552), .D(
        poly7_shifted[90]), .Z(n17240) );
  COND1XL U17248 ( .A(n17305), .B(n17471), .C(n17240), .Z(n10014) );
  CANR2X1 U17249 ( .A(n17453), .B(poly0_shifted[186]), .C(n17314), .D(
        poly0_shifted[204]), .Z(n17241) );
  COND1XL U17250 ( .A(n17316), .B(n17735), .C(n17241), .Z(n9391) );
  CANR2X1 U17251 ( .A(n18047), .B(poly0_shifted[154]), .C(n17671), .D(
        Poly0[154]), .Z(n17242) );
  COND1XL U17252 ( .A(n17674), .B(n17735), .C(n17242), .Z(n9423) );
  CANR2X1 U17253 ( .A(n18234), .B(poly0_shifted[58]), .C(n17500), .D(
        poly0_shifted[76]), .Z(n17243) );
  COND1XL U17254 ( .A(n17502), .B(n17305), .C(n17243), .Z(n9519) );
  CANR2X1 U17255 ( .A(n12625), .B(poly7_shifted[294]), .C(n16435), .D(
        poly7_shifted[282]), .Z(n17244) );
  COND1XL U17256 ( .A(n17305), .B(n12625), .C(n17244), .Z(n9822) );
  CANR2X1 U17257 ( .A(n15737), .B(poly3_shifted[40]), .C(n17245), .D(
        poly3_shifted[26]), .Z(n17246) );
  COND1XL U17258 ( .A(n17735), .B(n15737), .C(n17246), .Z(n8914) );
  CANR2X1 U17259 ( .A(n12598), .B(Poly12[58]), .C(n17714), .D(
        poly12_shifted[58]), .Z(n17247) );
  COND1XL U17260 ( .A(n17735), .B(n12598), .C(n17247), .Z(n10474) );
  CANR2X1 U17261 ( .A(n18018), .B(Poly7[26]), .C(n16644), .D(poly7_shifted[26]), .Z(n17248) );
  COND1XL U17262 ( .A(n17735), .B(n18018), .C(n17248), .Z(n10078) );
  CANR2X1 U17263 ( .A(n12211), .B(Poly2[26]), .C(n17508), .D(poly2_shifted[26]), .Z(n17249) );
  COND1XL U17264 ( .A(n17735), .B(n12211), .C(n17249), .Z(n8984) );
  CANR2XL U17265 ( .A(n18191), .B(poly1_shifted[293]), .C(n17640), .D(
        poly1_shifted[282]), .Z(n17250) );
  COND1XL U17266 ( .A(n17735), .B(n18191), .C(n17250), .Z(n9075) );
  CANR2X1 U17267 ( .A(n12299), .B(Poly1[58]), .C(n16312), .D(poly1_shifted[58]), .Z(n17251) );
  COND1XL U17268 ( .A(n17305), .B(n12299), .C(n17251), .Z(n9299) );
  CANR2X1 U17269 ( .A(n12401), .B(Poly7[410]), .C(n17449), .D(
        poly7_shifted[410]), .Z(n17252) );
  COND1XL U17270 ( .A(n17305), .B(n12401), .C(n17252), .Z(n9694) );
  CEOXL U17271 ( .A(Poly14[288]), .B(Poly14[294]), .Z(n17253) );
  CENX1 U17272 ( .A(Poly14[202]), .B(n17253), .Z(n17254) );
  CNR2XL U17273 ( .A(n17826), .B(n17254), .Z(n17255) );
  CANR1XL U17274 ( .A(poly14_shifted[234]), .B(n12202), .C(n17255), .Z(n17256)
         );
  COND1XL U17275 ( .A(n17735), .B(n12202), .C(n17256), .Z(n10187) );
  CANR2X1 U17276 ( .A(n12210), .B(poly1_shifted[197]), .C(n17466), .D(
        poly1_shifted[186]), .Z(n17257) );
  COND1XL U17277 ( .A(n17735), .B(n12210), .C(n17257), .Z(n9171) );
  CEOXL U17278 ( .A(Poly3[77]), .B(Poly3[83]), .Z(n17258) );
  CENX1 U17279 ( .A(Poly3[44]), .B(n17258), .Z(n17260) );
  CNR2XL U17280 ( .A(n17260), .B(n17259), .Z(n17261) );
  CANR1XL U17281 ( .A(Poly3[58]), .B(n17262), .C(n17261), .Z(n17263) );
  COND1XL U17282 ( .A(n17305), .B(n17589), .C(n17263), .Z(n8882) );
  CANR2X1 U17283 ( .A(n17982), .B(poly13_shifted[392]), .C(n17266), .D(
        poly13_shifted[378]), .Z(n17264) );
  COND1XL U17284 ( .A(n17735), .B(n17982), .C(n17264), .Z(n10682) );
  CANR2X1 U17285 ( .A(n17525), .B(poly14_shifted[74]), .C(n17613), .D(
        poly14_shifted[58]), .Z(n17265) );
  COND1XL U17286 ( .A(n17735), .B(n17525), .C(n17265), .Z(n10347) );
  CANR2X1 U17287 ( .A(n17969), .B(poly13_shifted[104]), .C(n17266), .D(
        poly13_shifted[90]), .Z(n17267) );
  COND1XL U17288 ( .A(n17735), .B(n17969), .C(n17267), .Z(n10970) );
  CANR2X1 U17289 ( .A(n18230), .B(Poly4[26]), .C(n17334), .D(poly4_shifted[26]), .Z(n17268) );
  COND1XL U17290 ( .A(n17735), .B(n18230), .C(n17268), .Z(n8830) );
  CANR2X1 U17291 ( .A(n12012), .B(poly1_shifted[101]), .C(n18234), .D(
        poly1_shifted[90]), .Z(n17269) );
  COND1XL U17292 ( .A(n17735), .B(n12012), .C(n17269), .Z(n9267) );
  CANR2XL U17293 ( .A(n18002), .B(poly14_shifted[42]), .C(poly14_shifted[26]), 
        .D(n18017), .Z(n17270) );
  COND1XL U17294 ( .A(n17305), .B(n18002), .C(n17270), .Z(n10379) );
  CANR2X1 U17295 ( .A(n17592), .B(Poly13[282]), .C(n17266), .D(
        poly13_shifted[282]), .Z(n17271) );
  COND1XL U17296 ( .A(n17305), .B(n17592), .C(n17271), .Z(n10778) );
  CANR2X1 U17297 ( .A(n17273), .B(poly7_shifted[230]), .C(n17545), .D(
        poly7_shifted[218]), .Z(n17272) );
  COND1XL U17298 ( .A(n17735), .B(n17273), .C(n17272), .Z(n9886) );
  CANR2X1 U17299 ( .A(n16425), .B(poly1_shifted[133]), .C(n17504), .D(
        poly1_shifted[122]), .Z(n17274) );
  COND1XL U17300 ( .A(n17305), .B(n16425), .C(n17274), .Z(n9235) );
  CANR2X1 U17301 ( .A(n12958), .B(poly14_shifted[106]), .C(n17965), .D(
        poly14_shifted[90]), .Z(n17275) );
  COND1XL U17302 ( .A(n17735), .B(n12958), .C(n17275), .Z(n10315) );
  CANR2X1 U17303 ( .A(n12932), .B(poly14_shifted[298]), .C(n17714), .D(
        poly14_shifted[282]), .Z(n17276) );
  COND1XL U17304 ( .A(n17735), .B(n12932), .C(n17276), .Z(n10123) );
  CANR2X1 U17305 ( .A(n17491), .B(poly13_shifted[520]), .C(n17508), .D(
        poly13_shifted[506]), .Z(n17277) );
  COND1XL U17306 ( .A(n17735), .B(n17491), .C(n17277), .Z(n10554) );
  CANR2X1 U17307 ( .A(n13124), .B(poly13_shifted[40]), .C(n17755), .D(
        poly13_shifted[26]), .Z(n17278) );
  COND1XL U17308 ( .A(n17305), .B(n13124), .C(n17278), .Z(n11034) );
  CANR2X1 U17309 ( .A(n16694), .B(poly14_shifted[266]), .C(n18234), .D(
        poly14_shifted[250]), .Z(n17279) );
  COND1XL U17310 ( .A(n17305), .B(n16694), .C(n17279), .Z(n10155) );
  CANR2X1 U17311 ( .A(n17974), .B(poly13_shifted[136]), .C(n17280), .D(
        poly13_shifted[122]), .Z(n17281) );
  COND1XL U17312 ( .A(n17735), .B(n17974), .C(n17281), .Z(n10938) );
  CANR2X1 U17313 ( .A(n13070), .B(poly7_shifted[166]), .C(n17334), .D(
        poly7_shifted[154]), .Z(n17282) );
  COND1XL U17314 ( .A(n17305), .B(n13070), .C(n17282), .Z(n9950) );
  CANR2X1 U17315 ( .A(n17987), .B(poly13_shifted[456]), .C(n17458), .D(
        poly13_shifted[442]), .Z(n17283) );
  COND1XL U17316 ( .A(n17735), .B(n17987), .C(n17283), .Z(n10618) );
  CANR2XL U17317 ( .A(n12009), .B(poly14_shifted[138]), .C(poly14_shifted[122]), .D(n18017), .Z(n17284) );
  COND1XL U17318 ( .A(n17735), .B(n12009), .C(n17284), .Z(n10283) );
  CANR2X1 U17319 ( .A(n17667), .B(poly13_shifted[232]), .C(n17285), .D(
        poly13_shifted[218]), .Z(n17286) );
  COND1XL U17320 ( .A(n17305), .B(n17667), .C(n17286), .Z(n10842) );
  CANR2X1 U17321 ( .A(n12997), .B(Poly12[26]), .C(n17552), .D(
        poly12_shifted[26]), .Z(n17287) );
  COND1XL U17322 ( .A(n17735), .B(n12997), .C(n17287), .Z(n10506) );
  CANR2X1 U17323 ( .A(n12977), .B(Poly7[186]), .C(n17288), .D(
        poly7_shifted[186]), .Z(n17289) );
  COND1XL U17324 ( .A(n17735), .B(n12977), .C(n17289), .Z(n9918) );
  CANR2X1 U17325 ( .A(n17217), .B(poly7_shifted[134]), .C(n17290), .D(
        poly7_shifted[122]), .Z(n17291) );
  COND1XL U17326 ( .A(n17735), .B(n17217), .C(n17291), .Z(n9982) );
  CANR2X1 U17327 ( .A(n18044), .B(Poly15[26]), .C(n17072), .D(
        poly15_shifted[26]), .Z(n17292) );
  COND1XL U17328 ( .A(n17735), .B(n18044), .C(n17292), .Z(n9611) );
  CANR2XL U17329 ( .A(n17332), .B(Poly1[346]), .C(n17285), .D(
        poly1_shifted[346]), .Z(n17293) );
  COND1XL U17330 ( .A(n17305), .B(n17332), .C(n17293), .Z(n9011) );
  CANR2X1 U17331 ( .A(n13014), .B(poly13_shifted[200]), .C(n17538), .D(
        poly13_shifted[186]), .Z(n17294) );
  COND1XL U17332 ( .A(n17305), .B(n13014), .C(n17294), .Z(n10874) );
  CANR2X1 U17333 ( .A(n13040), .B(poly7_shifted[358]), .C(n17295), .D(
        poly7_shifted[346]), .Z(n17296) );
  COND1XL U17334 ( .A(n17735), .B(n13040), .C(n17296), .Z(n9758) );
  CANR2X1 U17335 ( .A(n12900), .B(poly13_shifted[72]), .C(n17209), .D(
        poly13_shifted[58]), .Z(n17297) );
  COND1XL U17336 ( .A(n17735), .B(n12900), .C(n17297), .Z(n11002) );
  CANR2X1 U17337 ( .A(n17615), .B(poly13_shifted[328]), .C(n17298), .D(
        poly13_shifted[314]), .Z(n17299) );
  COND1XL U17338 ( .A(n17735), .B(n17615), .C(n17299), .Z(n10746) );
  CANR2X1 U17339 ( .A(n12008), .B(poly14_shifted[170]), .C(n16702), .D(
        poly14_shifted[154]), .Z(n17300) );
  COND1XL U17340 ( .A(n17735), .B(n12008), .C(n17300), .Z(n10251) );
  CANR2X1 U17341 ( .A(n18028), .B(poly7_shifted[326]), .C(n17266), .D(
        poly7_shifted[314]), .Z(n17301) );
  COND1XL U17342 ( .A(n17305), .B(n18028), .C(n17301), .Z(n9790) );
  CANR2X1 U17343 ( .A(n17595), .B(poly13_shifted[264]), .C(n17755), .D(
        poly13_shifted[250]), .Z(n17302) );
  COND1XL U17344 ( .A(n17735), .B(n17595), .C(n17302), .Z(n10810) );
  CANR2X1 U17345 ( .A(n17990), .B(poly13_shifted[488]), .C(n17640), .D(
        poly13_shifted[474]), .Z(n17303) );
  COND1XL U17346 ( .A(n17735), .B(n17990), .C(n17303), .Z(n10586) );
  CANR2X1 U17347 ( .A(n17603), .B(poly13_shifted[360]), .C(n17965), .D(
        poly13_shifted[346]), .Z(n17304) );
  COND1XL U17348 ( .A(n17305), .B(n17603), .C(n17304), .Z(n10714) );
  CND2XL U17349 ( .A(Poly2[65]), .B(Poly2[25]), .Z(n17311) );
  CNR2X1 U17350 ( .A(Poly2[65]), .B(Poly2[25]), .Z(n17312) );
  CNR2XL U17351 ( .A(n17307), .B(n17312), .Z(n17308) );
  CND2X1 U17352 ( .A(n17308), .B(n17311), .Z(n17309) );
  CANR2X1 U17353 ( .A(n17099), .B(poly0_shifted[165]), .C(n17314), .D(
        Poly0[165]), .Z(n17315) );
  COND1XL U17354 ( .A(n17316), .B(n11993), .C(n17315), .Z(n9412) );
  CANR2X1 U17355 ( .A(n17317), .B(Poly0[207]), .C(n17503), .D(Poly0[5]), .Z(
        n17318) );
  COND1XL U17356 ( .A(n17506), .B(n11991), .C(n17318), .Z(n9572) );
  CANR2XL U17357 ( .A(n13124), .B(poly13_shifted[19]), .C(n17607), .D(
        Poly13[519]), .Z(n17319) );
  COND1XL U17358 ( .A(n11987), .B(n13124), .C(n17319), .Z(n11055) );
  CANR2X1 U17359 ( .A(n17595), .B(poly13_shifted[243]), .C(n17613), .D(
        poly13_shifted[229]), .Z(n17320) );
  COND1XL U17360 ( .A(n11993), .B(n17595), .C(n17320), .Z(n10831) );
  CEOXL U17361 ( .A(Poly12[117]), .B(Poly12[21]), .Z(n17321) );
  CANR2X1 U17362 ( .A(n12598), .B(Poly12[37]), .C(n16502), .D(n17321), .Z(
        n17322) );
  COND1XL U17363 ( .A(n11985), .B(n12598), .C(n17322), .Z(n10495) );
  CANR2X1 U17364 ( .A(n17525), .B(poly14_shifted[53]), .C(n17401), .D(
        poly14_shifted[37]), .Z(n17323) );
  COND1XL U17365 ( .A(n11989), .B(n17525), .C(n17323), .Z(n10368) );
  CANR2X1 U17366 ( .A(n17987), .B(poly13_shifted[435]), .C(n17538), .D(
        poly13_shifted[421]), .Z(n17324) );
  COND1XL U17367 ( .A(n11983), .B(n17987), .C(n17324), .Z(n10639) );
  CANR2X1 U17368 ( .A(n17982), .B(poly13_shifted[371]), .C(poly13_shifted[357]), .D(n18017), .Z(n17325) );
  COND1XL U17369 ( .A(n11995), .B(n17982), .C(n17325), .Z(n10703) );
  CEOX1 U17370 ( .A(n17327), .B(n17326), .Z(n17372) );
  CENX1 U17371 ( .A(Poly4[22]), .B(n17328), .Z(n17329) );
  CENX1 U17372 ( .A(n17372), .B(n17329), .Z(n17331) );
  CMXI2X1 U17373 ( .A0(n18138), .A1(Poly4[39]), .S(n12153), .Z(n17330) );
  COND1XL U17374 ( .A(n17331), .B(n17959), .C(n17330), .Z(n8817) );
  CANR2XL U17375 ( .A(n17332), .B(Poly1[343]), .C(n17998), .D(
        poly1_shifted[343]), .Z(n17333) );
  COND1XL U17376 ( .A(n12000), .B(n17332), .C(n17333), .Z(n9014) );
  CANR2X1 U17377 ( .A(n18230), .B(Poly4[23]), .C(n17334), .D(poly4_shifted[23]), .Z(n17335) );
  COND1XL U17378 ( .A(n12000), .B(n18230), .C(n17335), .Z(n8833) );
  CANR2X1 U17379 ( .A(n17977), .B(poly13_shifted[165]), .C(n16702), .D(
        poly13_shifted[151]), .Z(n17336) );
  COND1XL U17380 ( .A(n12000), .B(n17977), .C(n17336), .Z(n10909) );
  CEOX1 U17381 ( .A(Poly3[41]), .B(Poly3[74]), .Z(n17337) );
  CENX1 U17382 ( .A(Poly3[80]), .B(n17337), .Z(n17338) );
  CNR2XL U17383 ( .A(n17959), .B(n17338), .Z(n17339) );
  CANR1XL U17384 ( .A(Poly3[55]), .B(n17587), .C(n17339), .Z(n17340) );
  COND1XL U17385 ( .A(n12000), .B(n17589), .C(n17340), .Z(n8885) );
  CIVXL U17386 ( .A(n17685), .Z(n17341) );
  CANR2X1 U17387 ( .A(n12211), .B(poly2_shifted[16]), .C(n16488), .D(n17341), 
        .Z(n17342) );
  COND1XL U17388 ( .A(n12005), .B(n12211), .C(n17342), .Z(n9006) );
  CANR2X1 U17389 ( .A(n17955), .B(poly9_shifted[79]), .C(n17343), .D(
        poly9_shifted[68]), .Z(n17344) );
  COND1XL U17390 ( .A(n12005), .B(n17955), .C(n17344), .Z(n11237) );
  CEOXL U17391 ( .A(Poly9[89]), .B(Poly9[110]), .Z(n17345) );
  CANR2X1 U17392 ( .A(n12262), .B(poly9_shifted[111]), .C(n17598), .D(n17345), 
        .Z(n17346) );
  COND1XL U17393 ( .A(n12005), .B(n12262), .C(n17346), .Z(n11205) );
  CANR2X1 U17394 ( .A(n17671), .B(Poly0[151]), .C(n17094), .D(
        poly0_shifted[151]), .Z(n17347) );
  COND1XL U17395 ( .A(n17674), .B(n12000), .C(n17347), .Z(n9426) );
  CANR2X1 U17396 ( .A(n17974), .B(poly13_shifted[133]), .C(n17348), .D(
        poly13_shifted[119]), .Z(n17349) );
  COND1XL U17397 ( .A(n12296), .B(n17974), .C(n17349), .Z(n10941) );
  CANR2X1 U17398 ( .A(n12012), .B(poly1_shifted[98]), .C(n17362), .D(
        poly1_shifted[87]), .Z(n17350) );
  COND1XL U17399 ( .A(n12296), .B(n12012), .C(n17350), .Z(n9270) );
  CANR2X1 U17400 ( .A(n13070), .B(poly7_shifted[163]), .C(n17705), .D(
        poly7_shifted[151]), .Z(n17351) );
  COND1XL U17401 ( .A(n12000), .B(n13070), .C(n17351), .Z(n9953) );
  CANR2X1 U17402 ( .A(n18044), .B(Poly15[23]), .C(n17352), .D(
        poly15_shifted[23]), .Z(n17353) );
  COND1XL U17403 ( .A(n12000), .B(n18044), .C(n17353), .Z(n9614) );
  CANR2X1 U17404 ( .A(n17332), .B(poly1_shifted[336]), .C(n17449), .D(
        poly1_shifted[325]), .Z(n17354) );
  COND1XL U17405 ( .A(n11981), .B(n17332), .C(n17354), .Z(n9032) );
  CANR2X1 U17406 ( .A(n12192), .B(Poly1[229]), .C(n17965), .D(
        poly1_shifted[229]), .Z(n17355) );
  COND1XL U17407 ( .A(n11989), .B(n12192), .C(n17355), .Z(n9128) );
  CANR2X1 U17408 ( .A(n15737), .B(poly3_shifted[19]), .C(n17356), .D(Poly3[75]), .Z(n17357) );
  COND1XL U17409 ( .A(n11989), .B(n15737), .C(n17357), .Z(n8935) );
  CANR2XL U17410 ( .A(n18234), .B(poly0_shifted[19]), .C(n17503), .D(Poly0[19]), .Z(n17358) );
  COND1XL U17411 ( .A(n17506), .B(n17661), .C(n17358), .Z(n9558) );
  CANR2X1 U17412 ( .A(n17552), .B(poly3_shifted[83]), .C(Poly3[83]), .D(n17359), .Z(n17360) );
  COND1XL U17413 ( .A(n17361), .B(n17661), .C(n17360), .Z(n8857) );
  CANR2X1 U17414 ( .A(n17362), .B(poly0_shifted[51]), .C(n17500), .D(
        poly0_shifted[69]), .Z(n17363) );
  COND1XL U17415 ( .A(n17502), .B(n17661), .C(n17363), .Z(n9526) );
  CMXI2X1 U17416 ( .A0(n17366), .A1(n17364), .S(Poly2[56]), .Z(n17365) );
  CND2IX1 U17417 ( .B(n17696), .A(n17365), .Z(n17369) );
  CND2X1 U17418 ( .A(n17366), .B(Poly2[56]), .Z(n17367) );
  COND1XL U17419 ( .A(n17368), .B(n17369), .C(n17367), .Z(n17370) );
  CMXI2XL U17420 ( .A0(n17370), .A1(n17369), .S(Poly2[68]), .Z(n17371) );
  COND1XL U17421 ( .A(n12005), .B(n17696), .C(n17371), .Z(n8942) );
  CEOX1 U17422 ( .A(Poly4[31]), .B(n17372), .Z(n17374) );
  CMXI2X1 U17423 ( .A0(n18167), .A1(Poly4[48]), .S(n12153), .Z(n17373) );
  COND1XL U17424 ( .A(n17374), .B(n17495), .C(n17373), .Z(n8808) );
  CANR2X1 U17425 ( .A(n17376), .B(Poly15[55]), .C(n17375), .D(
        poly15_shifted[55]), .Z(n17377) );
  COND1XL U17426 ( .A(n12000), .B(n17376), .C(n17377), .Z(n9582) );
  CANR2X1 U17427 ( .A(n17969), .B(poly13_shifted[82]), .C(n16919), .D(
        poly13_shifted[68]), .Z(n17378) );
  COND1XL U17428 ( .A(n17423), .B(n17969), .C(n17378), .Z(n10992) );
  CANR2X1 U17429 ( .A(n12008), .B(poly14_shifted[148]), .C(n16919), .D(
        poly14_shifted[132]), .Z(n17379) );
  COND1XL U17430 ( .A(n17442), .B(n12008), .C(n17379), .Z(n10273) );
  CANR2X1 U17431 ( .A(n13040), .B(poly7_shifted[336]), .C(n17535), .D(
        poly7_shifted[324]), .Z(n17380) );
  COND1XL U17432 ( .A(n17417), .B(n13040), .C(n17380), .Z(n9780) );
  CANR2X1 U17433 ( .A(n17977), .B(poly13_shifted[146]), .C(n17508), .D(
        poly13_shifted[132]), .Z(n17381) );
  COND1XL U17434 ( .A(n17423), .B(n17977), .C(n17381), .Z(n10928) );
  CANR2X1 U17435 ( .A(n15737), .B(poly3_shifted[18]), .C(n17094), .D(Poly3[74]), .Z(n17382) );
  COND1XL U17436 ( .A(n17442), .B(n15737), .C(n17382), .Z(n8936) );
  CIVX2 U17437 ( .A(n12004), .Z(n17417) );
  CANR2X1 U17438 ( .A(n12625), .B(poly7_shifted[272]), .C(n17383), .D(
        poly7_shifted[260]), .Z(n17384) );
  COND1XL U17439 ( .A(n17417), .B(n12625), .C(n17384), .Z(n9844) );
  CANR2X1 U17440 ( .A(n17603), .B(poly13_shifted[338]), .C(n17523), .D(
        poly13_shifted[324]), .Z(n17385) );
  COND1XL U17441 ( .A(n17423), .B(n17603), .C(n17385), .Z(n10736) );
  CANR2X1 U17442 ( .A(n17750), .B(Poly8[68]), .C(n17755), .D(poly8_shifted[68]), .Z(n17386) );
  COND1XL U17443 ( .A(n17442), .B(n17750), .C(n17386), .Z(n11333) );
  CEOXL U17444 ( .A(Poly14[300]), .B(Poly14[180]), .Z(n17387) );
  CANR2X1 U17445 ( .A(n12202), .B(Poly14[196]), .C(n17398), .D(n17387), .Z(
        n17388) );
  COND1XL U17446 ( .A(n17417), .B(n12202), .C(n17388), .Z(n10209) );
  CANR2X1 U17447 ( .A(n12932), .B(poly14_shifted[276]), .C(n17398), .D(
        poly14_shifted[260]), .Z(n17389) );
  COND1XL U17448 ( .A(n12005), .B(n12932), .C(n17389), .Z(n10145) );
  CANR2X1 U17449 ( .A(n12206), .B(poly7_shifted[368]), .C(n17390), .D(
        poly7_shifted[356]), .Z(n17391) );
  COND1XL U17450 ( .A(n17417), .B(n12206), .C(n17391), .Z(n9748) );
  CANR2X1 U17451 ( .A(n12401), .B(poly7_shifted[400]), .C(n17488), .D(
        poly7_shifted[388]), .Z(n17392) );
  COND1XL U17452 ( .A(n17417), .B(n12401), .C(n17392), .Z(n9716) );
  CEOXL U17453 ( .A(Poly14[298]), .B(Poly14[212]), .Z(n17393) );
  CANR2X1 U17454 ( .A(n16694), .B(poly14_shifted[244]), .C(n17285), .D(n17393), 
        .Z(n17394) );
  COND1XL U17455 ( .A(n12005), .B(n16694), .C(n17394), .Z(n10177) );
  CANR2X1 U17456 ( .A(n12287), .B(poly8_shifted[50]), .C(n16644), .D(
        poly8_shifted[36]), .Z(n17395) );
  COND1XL U17457 ( .A(n17417), .B(n12287), .C(n17395), .Z(n11365) );
  CANR2X1 U17458 ( .A(n17987), .B(poly13_shifted[434]), .C(n17401), .D(
        poly13_shifted[420]), .Z(n17396) );
  COND1XL U17459 ( .A(n12005), .B(n17987), .C(n17396), .Z(n10640) );
  CANR2X1 U17460 ( .A(n17217), .B(poly7_shifted[112]), .C(n17266), .D(
        poly7_shifted[100]), .Z(n17397) );
  COND1XL U17461 ( .A(n17417), .B(n17217), .C(n17397), .Z(n10004) );
  CANR2X1 U17462 ( .A(n13129), .B(poly14_shifted[180]), .C(n17398), .D(
        poly14_shifted[164]), .Z(n17399) );
  COND1XL U17463 ( .A(n17423), .B(n13129), .C(n17399), .Z(n10241) );
  CEOXL U17464 ( .A(Poly12[114]), .B(Poly12[84]), .Z(n17400) );
  CANR2X1 U17465 ( .A(n17652), .B(poly12_shifted[116]), .C(n17401), .D(n17400), 
        .Z(n17402) );
  COND1XL U17466 ( .A(n17423), .B(n17652), .C(n17402), .Z(n10432) );
  CANR2X1 U17467 ( .A(n18028), .B(poly7_shifted[304]), .C(n17655), .D(
        poly7_shifted[292]), .Z(n17403) );
  COND1XL U17468 ( .A(n17442), .B(n18028), .C(n17403), .Z(n9812) );
  CEOXL U17469 ( .A(Poly13[523]), .B(Poly13[278]), .Z(n17404) );
  CANR2X1 U17470 ( .A(n17615), .B(poly13_shifted[306]), .C(n17634), .D(n17404), 
        .Z(n17405) );
  COND1XL U17471 ( .A(n17423), .B(n17615), .C(n17405), .Z(n10768) );
  CANR2X1 U17472 ( .A(n17592), .B(poly13_shifted[274]), .C(n17560), .D(
        poly13_shifted[260]), .Z(n17406) );
  COND1XL U17473 ( .A(n17423), .B(n17592), .C(n17406), .Z(n10800) );
  CANR2X1 U17474 ( .A(n18002), .B(poly14_shifted[20]), .C(n17508), .D(
        Poly14[289]), .Z(n17407) );
  COND1XL U17475 ( .A(n17417), .B(n18002), .C(n17407), .Z(n10401) );
  CANR2X1 U17476 ( .A(n17525), .B(poly14_shifted[52]), .C(n17642), .D(
        poly14_shifted[36]), .Z(n17408) );
  COND1XL U17477 ( .A(n17423), .B(n17525), .C(n17408), .Z(n10369) );
  CEOXL U17478 ( .A(Poly10[40]), .B(Poly10[24]), .Z(n17409) );
  CANR2XL U17479 ( .A(n17411), .B(Poly10[36]), .C(n18234), .D(n17409), .Z(
        n17410) );
  COND1XL U17480 ( .A(n17442), .B(n17411), .C(n17410), .Z(n11067) );
  CANR2X1 U17481 ( .A(n17990), .B(poly13_shifted[466]), .C(n17755), .D(
        poly13_shifted[452]), .Z(n17412) );
  COND1XL U17482 ( .A(n17423), .B(n17990), .C(n17412), .Z(n10608) );
  CANR2X1 U17483 ( .A(n13070), .B(poly7_shifted[144]), .C(n17545), .D(
        poly7_shifted[132]), .Z(n17413) );
  COND1XL U17484 ( .A(n17442), .B(n13070), .C(n17413), .Z(n9972) );
  CANR2XL U17485 ( .A(n18191), .B(poly1_shifted[271]), .C(n17998), .D(
        poly1_shifted[260]), .Z(n17414) );
  COND1XL U17486 ( .A(n17417), .B(n18191), .C(n17414), .Z(n9097) );
  CANR2X1 U17487 ( .A(n17982), .B(poly13_shifted[370]), .C(n17538), .D(
        poly13_shifted[356]), .Z(n17415) );
  COND1XL U17488 ( .A(n17423), .B(n17982), .C(n17415), .Z(n10704) );
  CANR2X1 U17489 ( .A(n18018), .B(poly7_shifted[16]), .C(n17099), .D(
        Poly7[403]), .Z(n17416) );
  COND1XL U17490 ( .A(n17417), .B(n18018), .C(n17416), .Z(n10100) );
  CANR2X1 U17491 ( .A(n17491), .B(poly13_shifted[498]), .C(n16323), .D(
        poly13_shifted[484]), .Z(n17418) );
  COND1XL U17492 ( .A(n17442), .B(n17491), .C(n17418), .Z(n10576) );
  CANR2X1 U17493 ( .A(n16425), .B(poly1_shifted[111]), .C(n17099), .D(
        poly1_shifted[100]), .Z(n17419) );
  COND1XL U17494 ( .A(n17417), .B(n16425), .C(n17419), .Z(n9257) );
  CANR2X1 U17495 ( .A(n13014), .B(Poly13[164]), .C(n17466), .D(
        poly13_shifted[164]), .Z(n17420) );
  COND1XL U17496 ( .A(n17423), .B(n13014), .C(n17420), .Z(n10896) );
  CANR2XL U17497 ( .A(n12958), .B(poly14_shifted[84]), .C(n17634), .D(
        poly14_shifted[68]), .Z(n17421) );
  COND1XL U17498 ( .A(n17417), .B(n12958), .C(n17421), .Z(n10337) );
  CANR2X1 U17499 ( .A(n12900), .B(poly13_shifted[50]), .C(n17755), .D(
        poly13_shifted[36]), .Z(n17422) );
  COND1XL U17500 ( .A(n17423), .B(n12900), .C(n17422), .Z(n11024) );
  CANR2XL U17501 ( .A(n17610), .B(poly1_shifted[143]), .C(poly1_shifted[132]), 
        .D(n18017), .Z(n17424) );
  COND1XL U17502 ( .A(n12005), .B(n17610), .C(n17424), .Z(n9225) );
  CANR2X1 U17503 ( .A(n17667), .B(poly13_shifted[210]), .C(n17552), .D(
        poly13_shifted[196]), .Z(n17425) );
  COND1XL U17504 ( .A(n17442), .B(n17667), .C(n17425), .Z(n10864) );
  CANR2XL U17505 ( .A(n12009), .B(poly14_shifted[116]), .C(n18017), .D(
        poly14_shifted[100]), .Z(n17426) );
  COND1XL U17506 ( .A(n17423), .B(n12009), .C(n17426), .Z(n10305) );
  CANR2X1 U17507 ( .A(n17731), .B(poly9_shifted[15]), .C(n17449), .D(
        Poly9[109]), .Z(n17427) );
  COND1XL U17508 ( .A(n17442), .B(n17731), .C(n17427), .Z(n11301) );
  CANR2X1 U17509 ( .A(n12175), .B(Poly8[4]), .C(n17245), .D(Poly8[86]), .Z(
        n17428) );
  COND1XL U17510 ( .A(n17417), .B(n12175), .C(n17428), .Z(n11397) );
  CANR2X1 U17511 ( .A(n17430), .B(Poly13[516]), .C(n18234), .D(
        poly13_shifted[516]), .Z(n17429) );
  COND1XL U17512 ( .A(n17442), .B(n17430), .C(n17429), .Z(n10544) );
  CAN2XL U17513 ( .A(n18017), .B(Poly12[115]), .Z(n17431) );
  CANR1XL U17514 ( .A(poly12_shifted[20]), .B(n12997), .C(n17431), .Z(n17432)
         );
  COND1XL U17515 ( .A(n12005), .B(n12997), .C(n17432), .Z(n10528) );
  CENX1 U17516 ( .A(Poly12[111]), .B(Poly12[112]), .Z(n17433) );
  CENX1 U17517 ( .A(Poly12[52]), .B(n17433), .Z(n17434) );
  CANR2X1 U17518 ( .A(n12161), .B(poly12_shifted[84]), .C(n17705), .D(n17434), 
        .Z(n17435) );
  COND1XL U17519 ( .A(n12005), .B(n12161), .C(n17435), .Z(n10464) );
  CANR2X1 U17520 ( .A(n17053), .B(poly1_shifted[207]), .C(n16479), .D(
        poly1_shifted[196]), .Z(n17436) );
  COND1XL U17521 ( .A(n12005), .B(n17053), .C(n17436), .Z(n9161) );
  CANR2X1 U17522 ( .A(n17595), .B(poly13_shifted[242]), .C(n17755), .D(
        poly13_shifted[228]), .Z(n17437) );
  COND1XL U17523 ( .A(n17442), .B(n17595), .C(n17437), .Z(n10832) );
  CEOXL U17524 ( .A(Poly9[114]), .B(Poly9[25]), .Z(n17438) );
  CANR2X1 U17525 ( .A(n13351), .B(poly9_shifted[47]), .C(n17538), .D(n17438), 
        .Z(n17439) );
  COND1XL U17526 ( .A(n17442), .B(n13351), .C(n17439), .Z(n11269) );
  CANR2X1 U17527 ( .A(n17574), .B(poly7_shifted[240]), .C(n17535), .D(
        poly7_shifted[228]), .Z(n17440) );
  COND1XL U17528 ( .A(n17423), .B(n17574), .C(n17440), .Z(n9876) );
  CANR2X1 U17529 ( .A(n17974), .B(poly13_shifted[114]), .C(n17705), .D(
        poly13_shifted[100]), .Z(n17441) );
  COND1XL U17530 ( .A(n17442), .B(n17974), .C(n17441), .Z(n10960) );
  CANR2XL U17531 ( .A(n17444), .B(Poly14[292]), .C(n17998), .D(
        poly14_shifted[292]), .Z(n17443) );
  COND1XL U17532 ( .A(n12005), .B(n17444), .C(n17443), .Z(n10113) );
  CANR2X1 U17533 ( .A(n18018), .B(Poly7[23]), .C(n17655), .D(poly7_shifted[23]), .Z(n17445) );
  COND1XL U17534 ( .A(n12296), .B(n18018), .C(n17445), .Z(n10081) );
  CANR2X1 U17535 ( .A(n12008), .B(poly14_shifted[167]), .C(n17072), .D(
        poly14_shifted[151]), .Z(n17446) );
  COND1XL U17536 ( .A(n12296), .B(n12008), .C(n17446), .Z(n10254) );
  CANR2X1 U17537 ( .A(n17273), .B(poly7_shifted[227]), .C(n17535), .D(
        poly7_shifted[215]), .Z(n17447) );
  COND1XL U17538 ( .A(n12296), .B(n17273), .C(n17447), .Z(n9889) );
  CANR2X1 U17539 ( .A(n17969), .B(poly13_shifted[101]), .C(n17144), .D(
        poly13_shifted[87]), .Z(n17448) );
  COND1XL U17540 ( .A(n12000), .B(n17969), .C(n17448), .Z(n10973) );
  CANR2X1 U17541 ( .A(n17610), .B(Poly1[151]), .C(n17449), .D(
        poly1_shifted[151]), .Z(n17450) );
  COND1XL U17542 ( .A(n12000), .B(n17610), .C(n17450), .Z(n9206) );
  CANR2X1 U17543 ( .A(n17525), .B(poly14_shifted[71]), .C(n17063), .D(
        poly14_shifted[55]), .Z(n17451) );
  COND1XL U17544 ( .A(n12000), .B(n17525), .C(n17451), .Z(n10350) );
  CANR2X1 U17545 ( .A(n12997), .B(Poly12[23]), .C(n17613), .D(
        poly12_shifted[23]), .Z(n17452) );
  COND1XL U17546 ( .A(n12296), .B(n12997), .C(n17452), .Z(n10509) );
  CANR2X1 U17547 ( .A(n13040), .B(poly7_shifted[355]), .C(n17453), .D(
        poly7_shifted[343]), .Z(n17454) );
  COND1XL U17548 ( .A(n12296), .B(n13040), .C(n17454), .Z(n9761) );
  CANR2XL U17549 ( .A(n12958), .B(poly14_shifted[103]), .C(n17238), .D(
        poly14_shifted[87]), .Z(n17455) );
  COND1XL U17550 ( .A(n12296), .B(n12958), .C(n17455), .Z(n10318) );
  CANR2X1 U17551 ( .A(n12211), .B(Poly2[23]), .C(n16985), .D(poly2_shifted[23]), .Z(n17456) );
  COND1XL U17552 ( .A(n12000), .B(n12211), .C(n17456), .Z(n8987) );
  CANR2X1 U17553 ( .A(n17667), .B(poly13_shifted[229]), .C(n17508), .D(
        poly13_shifted[215]), .Z(n17457) );
  COND1XL U17554 ( .A(n12000), .B(n17667), .C(n17457), .Z(n10845) );
  CANR2X1 U17555 ( .A(n12977), .B(Poly7[183]), .C(n17458), .D(
        poly7_shifted[183]), .Z(n17459) );
  COND1XL U17556 ( .A(n12296), .B(n12977), .C(n17459), .Z(n9921) );
  CANR2X1 U17557 ( .A(n12009), .B(poly14_shifted[135]), .C(n17063), .D(
        poly14_shifted[119]), .Z(n17460) );
  COND1XL U17558 ( .A(n12296), .B(n12009), .C(n17460), .Z(n10286) );
  CANR2X1 U17559 ( .A(n17217), .B(poly7_shifted[131]), .C(n17535), .D(
        poly7_shifted[119]), .Z(n17461) );
  COND1XL U17560 ( .A(n12296), .B(n17217), .C(n17461), .Z(n9985) );
  CANR2X1 U17561 ( .A(n17982), .B(poly13_shifted[389]), .C(n17755), .D(
        poly13_shifted[375]), .Z(n17462) );
  COND1XL U17562 ( .A(n12296), .B(n17982), .C(n17462), .Z(n10685) );
  CANR2X1 U17563 ( .A(n16425), .B(poly1_shifted[130]), .C(n17642), .D(
        poly1_shifted[119]), .Z(n17463) );
  COND1XL U17564 ( .A(n12000), .B(n16425), .C(n17463), .Z(n9238) );
  CANR2X1 U17565 ( .A(n17592), .B(Poly13[279]), .C(n17401), .D(
        poly13_shifted[279]), .Z(n17464) );
  COND1XL U17566 ( .A(n12296), .B(n17592), .C(n17464), .Z(n10781) );
  CANR2X1 U17567 ( .A(n12401), .B(Poly7[407]), .C(n16307), .D(
        poly7_shifted[407]), .Z(n17465) );
  COND1XL U17568 ( .A(n12000), .B(n12401), .C(n17465), .Z(n9697) );
  CANR2X1 U17569 ( .A(n17987), .B(poly13_shifted[453]), .C(n17466), .D(
        poly13_shifted[439]), .Z(n17467) );
  COND1XL U17570 ( .A(n12296), .B(n17987), .C(n17467), .Z(n10621) );
  CANR2X1 U17571 ( .A(n18002), .B(poly14_shifted[39]), .C(n17449), .D(
        poly14_shifted[23]), .Z(n17468) );
  COND1XL U17572 ( .A(n12000), .B(n18002), .C(n17468), .Z(n10382) );
  CANR2X1 U17573 ( .A(n12625), .B(poly7_shifted[291]), .C(n17705), .D(
        poly7_shifted[279]), .Z(n17469) );
  COND1XL U17574 ( .A(n12296), .B(n12625), .C(n17469), .Z(n9825) );
  CANR2X1 U17575 ( .A(n17471), .B(poly7_shifted[99]), .C(n17552), .D(
        poly7_shifted[87]), .Z(n17470) );
  COND1XL U17576 ( .A(n12296), .B(n17471), .C(n17470), .Z(n10017) );
  CANR2X1 U17577 ( .A(n12161), .B(Poly12[87]), .C(n18234), .D(
        poly12_shifted[87]), .Z(n17472) );
  COND1XL U17578 ( .A(n12296), .B(n12161), .C(n17472), .Z(n10445) );
  CANR2X1 U17579 ( .A(n12932), .B(poly14_shifted[295]), .C(n18234), .D(
        poly14_shifted[279]), .Z(n17473) );
  COND1XL U17580 ( .A(n12296), .B(n12932), .C(n17473), .Z(n10126) );
  CANR2X1 U17581 ( .A(n12206), .B(poly7_shifted[387]), .C(n17362), .D(
        poly7_shifted[375]), .Z(n17474) );
  COND1XL U17582 ( .A(n12296), .B(n12206), .C(n17474), .Z(n9729) );
  CANR2X1 U17583 ( .A(n18191), .B(poly1_shifted[290]), .C(n18047), .D(
        poly1_shifted[279]), .Z(n17475) );
  COND1XL U17584 ( .A(n12000), .B(n18191), .C(n17475), .Z(n9078) );
  CANR2X1 U17585 ( .A(n12900), .B(poly13_shifted[69]), .C(n16323), .D(
        poly13_shifted[55]), .Z(n17476) );
  COND1XL U17586 ( .A(n12296), .B(n12900), .C(n17476), .Z(n11005) );
  CANR2X1 U17587 ( .A(n17595), .B(poly13_shifted[261]), .C(n17755), .D(
        poly13_shifted[247]), .Z(n17477) );
  COND1XL U17588 ( .A(n12296), .B(n17595), .C(n17477), .Z(n10813) );
  CEOXL U17589 ( .A(Poly14[285]), .B(Poly14[291]), .Z(n17478) );
  CENX1 U17590 ( .A(Poly14[199]), .B(n17478), .Z(n17479) );
  CNR2XL U17591 ( .A(n17479), .B(n17826), .Z(n17480) );
  CANR1XL U17592 ( .A(poly14_shifted[231]), .B(n12202), .C(n17480), .Z(n17481)
         );
  COND1XL U17593 ( .A(n12296), .B(n12202), .C(n17481), .Z(n10190) );
  CANR2X1 U17594 ( .A(n17990), .B(poly13_shifted[485]), .C(n17266), .D(
        poly13_shifted[471]), .Z(n17482) );
  COND1XL U17595 ( .A(n12000), .B(n17990), .C(n17482), .Z(n10589) );
  CANR2X1 U17596 ( .A(n13124), .B(poly13_shifted[37]), .C(n17668), .D(
        poly13_shifted[23]), .Z(n17483) );
  COND1XL U17597 ( .A(n12296), .B(n13124), .C(n17483), .Z(n11037) );
  CANR2X1 U17598 ( .A(n18198), .B(poly1_shifted[322]), .C(n17552), .D(
        poly1_shifted[311]), .Z(n17484) );
  COND1XL U17599 ( .A(n12000), .B(n18198), .C(n17484), .Z(n9046) );
  CANR2XL U17600 ( .A(n17603), .B(poly13_shifted[357]), .C(poly13_shifted[343]), .D(n18017), .Z(n17485) );
  COND1XL U17601 ( .A(n12296), .B(n17603), .C(n17485), .Z(n10717) );
  CANR2X1 U17602 ( .A(n16694), .B(poly14_shifted[263]), .C(n17965), .D(
        poly14_shifted[247]), .Z(n17486) );
  COND1XL U17603 ( .A(n12296), .B(n16694), .C(n17486), .Z(n10158) );
  CANR2XL U17604 ( .A(n12598), .B(Poly12[55]), .C(n18017), .D(
        poly12_shifted[55]), .Z(n17487) );
  COND1XL U17605 ( .A(n12296), .B(n12598), .C(n17487), .Z(n10477) );
  CANR2X1 U17606 ( .A(n17615), .B(poly13_shifted[325]), .C(n17488), .D(
        poly13_shifted[311]), .Z(n17489) );
  COND1XL U17607 ( .A(n12000), .B(n17615), .C(n17489), .Z(n10749) );
  CANR2X1 U17608 ( .A(n17731), .B(Poly9[23]), .C(n17705), .D(poly9_shifted[23]), .Z(n17490) );
  COND1XL U17609 ( .A(n12000), .B(n17731), .C(n17490), .Z(n11282) );
  CANR2XL U17610 ( .A(n17491), .B(poly13_shifted[517]), .C(n17285), .D(
        poly13_shifted[503]), .Z(n17492) );
  COND1XL U17611 ( .A(n12000), .B(n17491), .C(n17492), .Z(n10557) );
  CANR2X1 U17612 ( .A(n18028), .B(poly7_shifted[323]), .C(n17655), .D(
        poly7_shifted[311]), .Z(n17493) );
  COND1XL U17613 ( .A(n12296), .B(n18028), .C(n17493), .Z(n9793) );
  CEOXL U17614 ( .A(Poly12[125]), .B(Poly12[126]), .Z(n17494) );
  CENX1 U17615 ( .A(Poly12[66]), .B(n17494), .Z(n17496) );
  CNR2XL U17616 ( .A(n17496), .B(n17495), .Z(n17497) );
  CANR1XL U17617 ( .A(Poly12[82]), .B(n12161), .C(n17497), .Z(n17498) );
  COND1XL U17618 ( .A(n17549), .B(n12161), .C(n17498), .Z(n10450) );
  CANR2X1 U17619 ( .A(n16695), .B(poly0_shifted[146]), .C(poly0_shifted[164]), 
        .D(n17671), .Z(n17499) );
  COND1XL U17620 ( .A(n17674), .B(n17549), .C(n17499), .Z(n9431) );
  CANR2X1 U17621 ( .A(n17705), .B(poly0_shifted[50]), .C(poly0_shifted[68]), 
        .D(n17500), .Z(n17501) );
  COND1XL U17622 ( .A(n17502), .B(n17549), .C(n17501), .Z(n9527) );
  CANR2X1 U17623 ( .A(n17504), .B(poly0_shifted[18]), .C(n17503), .D(Poly0[18]), .Z(n17505) );
  COND1XL U17624 ( .A(n17506), .B(n17549), .C(n17505), .Z(n9559) );
  CIVX2 U17625 ( .A(n18210), .Z(n17571) );
  CANR2X1 U17626 ( .A(n17987), .B(poly13_shifted[448]), .C(n17063), .D(
        poly13_shifted[434]), .Z(n17507) );
  COND1XL U17627 ( .A(n17571), .B(n17987), .C(n17507), .Z(n10626) );
  CIVX2 U17628 ( .A(n18210), .Z(n17558) );
  CANR2X1 U17629 ( .A(n17977), .B(poly13_shifted[160]), .C(n17508), .D(
        poly13_shifted[146]), .Z(n17509) );
  COND1XL U17630 ( .A(n17558), .B(n17977), .C(n17509), .Z(n10914) );
  CIVX2 U17631 ( .A(n18210), .Z(n17569) );
  CANR2X1 U17632 ( .A(n12211), .B(Poly2[18]), .C(n17209), .D(poly2_shifted[18]), .Z(n17510) );
  COND1XL U17633 ( .A(n17569), .B(n12211), .C(n17510), .Z(n8992) );
  CANR2X1 U17634 ( .A(n17610), .B(poly1_shifted[157]), .C(n17598), .D(
        poly1_shifted[146]), .Z(n17511) );
  COND1XL U17635 ( .A(n17567), .B(n17610), .C(n17511), .Z(n9211) );
  CIVX2 U17636 ( .A(n18210), .Z(n17551) );
  CANR2X1 U17637 ( .A(n18002), .B(poly14_shifted[34]), .C(n17523), .D(
        poly14_shifted[18]), .Z(n17512) );
  COND1XL U17638 ( .A(n17551), .B(n18002), .C(n17512), .Z(n10387) );
  CANR2X1 U17639 ( .A(n17955), .B(poly9_shifted[93]), .C(n16702), .D(
        poly9_shifted[82]), .Z(n17513) );
  COND1XL U17640 ( .A(n17571), .B(n17955), .C(n17513), .Z(n11223) );
  CANR2X1 U17641 ( .A(n17273), .B(poly7_shifted[222]), .C(n16427), .D(
        poly7_shifted[210]), .Z(n17514) );
  COND1XL U17642 ( .A(n17571), .B(n17273), .C(n17514), .Z(n9894) );
  CANR2X1 U17643 ( .A(n12958), .B(poly14_shifted[98]), .C(n17527), .D(
        poly14_shifted[82]), .Z(n17515) );
  COND1XL U17644 ( .A(n17549), .B(n12958), .C(n17515), .Z(n10323) );
  CANR2X1 U17645 ( .A(n12401), .B(Poly7[402]), .C(n17552), .D(
        poly7_shifted[402]), .Z(n17516) );
  COND1XL U17646 ( .A(n17569), .B(n12401), .C(n17516), .Z(n9702) );
  CANR2X1 U17647 ( .A(n13040), .B(poly7_shifted[350]), .C(n17280), .D(
        poly7_shifted[338]), .Z(n17517) );
  COND1XL U17648 ( .A(n17549), .B(n13040), .C(n17517), .Z(n9766) );
  CANR2X1 U17649 ( .A(n18028), .B(poly7_shifted[318]), .C(n17527), .D(
        poly7_shifted[306]), .Z(n17518) );
  COND1XL U17650 ( .A(n17549), .B(n18028), .C(n17518), .Z(n9798) );
  CANR2X1 U17651 ( .A(n18230), .B(Poly4[18]), .C(n17552), .D(poly4_shifted[18]), .Z(n17519) );
  COND1XL U17652 ( .A(n17569), .B(n18230), .C(n17519), .Z(n8838) );
  CANR2X1 U17653 ( .A(n15737), .B(poly3_shifted[32]), .C(n17504), .D(
        poly3_shifted[18]), .Z(n17520) );
  COND1XL U17654 ( .A(n17567), .B(n15737), .C(n17520), .Z(n8922) );
  CANR2X1 U17655 ( .A(n17667), .B(poly13_shifted[224]), .C(n17538), .D(
        poly13_shifted[210]), .Z(n17521) );
  COND1XL U17656 ( .A(n17571), .B(n17667), .C(n17521), .Z(n10850) );
  CANR2X1 U17657 ( .A(n17652), .B(Poly12[114]), .C(n17655), .D(
        poly12_shifted[114]), .Z(n17522) );
  COND1XL U17658 ( .A(n17551), .B(n17652), .C(n17522), .Z(n10418) );
  CANR2X1 U17659 ( .A(n17525), .B(poly14_shifted[66]), .C(n17523), .D(
        poly14_shifted[50]), .Z(n17524) );
  COND1XL U17660 ( .A(n17551), .B(n17525), .C(n17524), .Z(n10355) );
  CANR2X1 U17661 ( .A(n17603), .B(poly13_shifted[352]), .C(n17362), .D(
        poly13_shifted[338]), .Z(n17526) );
  COND1XL U17662 ( .A(n17569), .B(n17603), .C(n17526), .Z(n10722) );
  CANR2X1 U17663 ( .A(n12009), .B(poly14_shifted[130]), .C(n17527), .D(
        poly14_shifted[114]), .Z(n17528) );
  COND1XL U17664 ( .A(n17549), .B(n12009), .C(n17528), .Z(n10291) );
  CANR2X1 U17665 ( .A(n13351), .B(poly9_shifted[61]), .C(n18234), .D(
        poly9_shifted[50]), .Z(n17529) );
  COND1XL U17666 ( .A(n17571), .B(n13351), .C(n17529), .Z(n11255) );
  CANR2X1 U17667 ( .A(n17969), .B(poly13_shifted[96]), .C(n17348), .D(
        poly13_shifted[82]), .Z(n17530) );
  COND1XL U17668 ( .A(n17551), .B(n17969), .C(n17530), .Z(n10978) );
  CANR2X1 U17669 ( .A(n17491), .B(poly13_shifted[512]), .C(n18234), .D(
        poly13_shifted[498]), .Z(n17531) );
  COND1XL U17670 ( .A(n17551), .B(n17491), .C(n17531), .Z(n10562) );
  CANR2X1 U17671 ( .A(n17974), .B(poly13_shifted[128]), .C(n17545), .D(
        poly13_shifted[114]), .Z(n17532) );
  COND1XL U17672 ( .A(n17551), .B(n17974), .C(n17532), .Z(n10946) );
  CANR2X1 U17673 ( .A(n17471), .B(poly7_shifted[94]), .C(n17533), .D(
        poly7_shifted[82]), .Z(n17534) );
  COND1XL U17674 ( .A(n17571), .B(n17471), .C(n17534), .Z(n10022) );
  CANR2X1 U17675 ( .A(n17574), .B(Poly7[242]), .C(n17535), .D(
        poly7_shifted[242]), .Z(n17536) );
  COND1XL U17676 ( .A(n17571), .B(n17574), .C(n17536), .Z(n9862) );
  CANR2X1 U17677 ( .A(n12997), .B(Poly12[18]), .C(n17755), .D(
        poly12_shifted[18]), .Z(n17537) );
  COND1XL U17678 ( .A(n17551), .B(n12997), .C(n17537), .Z(n10514) );
  CANR2X1 U17679 ( .A(n17982), .B(poly13_shifted[384]), .C(n17538), .D(
        poly13_shifted[370]), .Z(n17539) );
  COND1XL U17680 ( .A(n17558), .B(n17982), .C(n17539), .Z(n10690) );
  CANR2X1 U17681 ( .A(n12900), .B(poly13_shifted[64]), .C(n17755), .D(
        poly13_shifted[50]), .Z(n17540) );
  COND1XL U17682 ( .A(n17558), .B(n12900), .C(n17540), .Z(n11010) );
  CANR2X1 U17683 ( .A(n12625), .B(poly7_shifted[286]), .C(n17642), .D(
        poly7_shifted[274]), .Z(n17541) );
  COND1XL U17684 ( .A(n17569), .B(n12625), .C(n17541), .Z(n9830) );
  CANR2X1 U17685 ( .A(n12932), .B(poly14_shifted[290]), .C(n17508), .D(
        poly14_shifted[274]), .Z(n17542) );
  COND1XL U17686 ( .A(n17551), .B(n12932), .C(n17542), .Z(n10131) );
  CANR2X1 U17687 ( .A(n12012), .B(poly1_shifted[93]), .C(n17383), .D(
        poly1_shifted[82]), .Z(n17543) );
  COND1XL U17688 ( .A(n17567), .B(n12012), .C(n17543), .Z(n9275) );
  CANR2XL U17689 ( .A(n17592), .B(Poly13[274]), .C(n17607), .D(
        poly13_shifted[274]), .Z(n17544) );
  COND1XL U17690 ( .A(n17558), .B(n17592), .C(n17544), .Z(n10786) );
  CANR2X1 U17691 ( .A(n13124), .B(poly13_shifted[32]), .C(n17545), .D(
        poly13_shifted[18]), .Z(n17546) );
  COND1XL U17692 ( .A(n17551), .B(n13124), .C(n17546), .Z(n11042) );
  CANR2XL U17693 ( .A(n18191), .B(poly1_shifted[285]), .C(n17634), .D(
        poly1_shifted[274]), .Z(n17547) );
  COND1XL U17694 ( .A(n17567), .B(n18191), .C(n17547), .Z(n9083) );
  CANR2X1 U17695 ( .A(n12008), .B(poly14_shifted[162]), .C(n16435), .D(
        poly14_shifted[146]), .Z(n17548) );
  COND1XL U17696 ( .A(n17549), .B(n12008), .C(n17548), .Z(n10259) );
  CANR2X1 U17697 ( .A(n17595), .B(poly13_shifted[256]), .C(n17552), .D(
        poly13_shifted[242]), .Z(n17550) );
  COND1XL U17698 ( .A(n17551), .B(n17595), .C(n17550), .Z(n10818) );
  CANR2X1 U17699 ( .A(n13070), .B(poly7_shifted[158]), .C(n17552), .D(
        poly7_shifted[146]), .Z(n17553) );
  COND1XL U17700 ( .A(n17569), .B(n13070), .C(n17553), .Z(n9958) );
  CANR2X1 U17701 ( .A(n12977), .B(Poly7[178]), .C(n17655), .D(
        poly7_shifted[178]), .Z(n17554) );
  COND1XL U17702 ( .A(n17567), .B(n12977), .C(n17554), .Z(n9926) );
  CANR2XL U17703 ( .A(n16425), .B(poly1_shifted[125]), .C(poly1_shifted[114]), 
        .D(n18017), .Z(n17555) );
  COND1XL U17704 ( .A(n17567), .B(n16425), .C(n17555), .Z(n9243) );
  CANR2X1 U17705 ( .A(n12185), .B(Poly11[18]), .C(n17453), .D(
        poly11_shifted[18]), .Z(n17556) );
  COND1XL U17706 ( .A(n17571), .B(n12185), .C(n17556), .Z(n11171) );
  CANR2X1 U17707 ( .A(n17615), .B(poly13_shifted[320]), .C(n17634), .D(
        poly13_shifted[306]), .Z(n17557) );
  COND1XL U17708 ( .A(n17558), .B(n17615), .C(n17557), .Z(n10754) );
  CANR2X1 U17709 ( .A(n17990), .B(poly13_shifted[480]), .C(n17755), .D(
        poly13_shifted[466]), .Z(n17559) );
  COND1XL U17710 ( .A(n17569), .B(n17990), .C(n17559), .Z(n10594) );
  CANR2X1 U17711 ( .A(n17332), .B(Poly1[338]), .C(n17560), .D(
        poly1_shifted[338]), .Z(n17561) );
  COND1XL U17712 ( .A(n17569), .B(n17332), .C(n17561), .Z(n9019) );
  CANR2X1 U17713 ( .A(n12206), .B(poly7_shifted[382]), .C(n16372), .D(
        poly7_shifted[370]), .Z(n17562) );
  COND1XL U17714 ( .A(n17569), .B(n12206), .C(n17562), .Z(n9734) );
  CANR2X1 U17715 ( .A(n18018), .B(poly7_shifted[30]), .C(n17523), .D(
        poly7_shifted[18]), .Z(n17563) );
  COND1XL U17716 ( .A(n17571), .B(n17564), .C(n17563), .Z(n10086) );
  CANR2X1 U17717 ( .A(n12210), .B(poly1_shifted[189]), .C(n16307), .D(
        poly1_shifted[178]), .Z(n17565) );
  COND1XL U17718 ( .A(n17567), .B(n12210), .C(n17565), .Z(n9179) );
  CANR2X1 U17719 ( .A(n18044), .B(Poly15[18]), .C(n18047), .D(
        poly15_shifted[18]), .Z(n17566) );
  COND1XL U17720 ( .A(n17567), .B(n18044), .C(n17566), .Z(n9619) );
  CANR2X1 U17721 ( .A(n12170), .B(Poly7[50]), .C(n17598), .D(poly7_shifted[50]), .Z(n17568) );
  COND1XL U17722 ( .A(n17569), .B(n12170), .C(n17568), .Z(n10054) );
  CANR2X1 U17723 ( .A(n17217), .B(poly7_shifted[126]), .C(n17105), .D(
        poly7_shifted[114]), .Z(n17570) );
  COND1XL U17724 ( .A(n17571), .B(n17217), .C(n17570), .Z(n9990) );
  CANR2XL U17725 ( .A(n18044), .B(Poly15[19]), .C(poly15_shifted[19]), .D(
        n18017), .Z(n17572) );
  COND1XL U17726 ( .A(n17658), .B(n18044), .C(n17572), .Z(n9618) );
  CANR2XL U17727 ( .A(n17574), .B(Poly7[243]), .C(poly7_shifted[243]), .D(
        n18017), .Z(n17573) );
  COND1XL U17728 ( .A(n17664), .B(n17574), .C(n17573), .Z(n9861) );
  CANR2X1 U17729 ( .A(n17273), .B(poly7_shifted[223]), .C(n18234), .D(
        poly7_shifted[211]), .Z(n17575) );
  COND1XL U17730 ( .A(n17658), .B(n17273), .C(n17575), .Z(n9893) );
  CANR2X1 U17731 ( .A(n17376), .B(Poly15[51]), .C(n17523), .D(
        poly15_shifted[51]), .Z(n17576) );
  COND1XL U17732 ( .A(n17664), .B(n17376), .C(n17576), .Z(n9586) );
  CANR2X1 U17733 ( .A(n15737), .B(poly3_shifted[33]), .C(n16435), .D(
        poly3_shifted[19]), .Z(n17577) );
  COND1XL U17734 ( .A(n17673), .B(n15737), .C(n17577), .Z(n8921) );
  CANR2X1 U17735 ( .A(n12210), .B(poly1_shifted[190]), .C(n17121), .D(
        poly1_shifted[179]), .Z(n17578) );
  COND1XL U17736 ( .A(n17673), .B(n12210), .C(n17578), .Z(n9178) );
  CENX1 U17737 ( .A(Poly4[34]), .B(Poly4[59]), .Z(n17579) );
  CENX1 U17738 ( .A(n17580), .B(n17579), .Z(n17581) );
  CNR2XL U17739 ( .A(n17581), .B(n17826), .Z(n17582) );
  CANR1XL U17740 ( .A(Poly4[51]), .B(n12153), .C(n17582), .Z(n17583) );
  COND1XL U17741 ( .A(n17673), .B(n12153), .C(n17583), .Z(n8805) );
  CEOXL U17742 ( .A(Poly3[70]), .B(Poly3[76]), .Z(n17584) );
  CENX1 U17743 ( .A(Poly3[37]), .B(n17584), .Z(n17585) );
  CNR2XL U17744 ( .A(n17829), .B(n17585), .Z(n17586) );
  CANR1XL U17745 ( .A(Poly3[51]), .B(n17587), .C(n17586), .Z(n17588) );
  COND1XL U17746 ( .A(n17673), .B(n17589), .C(n17588), .Z(n8889) );
  CIVX2 U17747 ( .A(n18176), .Z(n17664) );
  CANR2X1 U17748 ( .A(n13129), .B(Poly14[179]), .C(n16427), .D(
        poly14_shifted[179]), .Z(n17590) );
  COND1XL U17749 ( .A(n17664), .B(n13129), .C(n17590), .Z(n10226) );
  CANR2X1 U17750 ( .A(n17592), .B(Poly13[275]), .C(n17755), .D(
        poly13_shifted[275]), .Z(n17591) );
  COND1XL U17751 ( .A(n17664), .B(n17592), .C(n17591), .Z(n10785) );
  CANR2X1 U17752 ( .A(n12932), .B(poly14_shifted[291]), .C(n17714), .D(
        poly14_shifted[275]), .Z(n17593) );
  COND1XL U17753 ( .A(n17664), .B(n12932), .C(n17593), .Z(n10130) );
  CIVX2 U17754 ( .A(n18176), .Z(n17658) );
  CANR2X1 U17755 ( .A(n17595), .B(poly13_shifted[257]), .C(n17449), .D(
        poly13_shifted[243]), .Z(n17594) );
  COND1XL U17756 ( .A(n17658), .B(n17595), .C(n17594), .Z(n10817) );
  CANR2X1 U17757 ( .A(n12401), .B(Poly7[403]), .C(n16488), .D(
        poly7_shifted[403]), .Z(n17596) );
  COND1XL U17758 ( .A(n17664), .B(n12401), .C(n17596), .Z(n9701) );
  CANR2X1 U17759 ( .A(n12170), .B(Poly7[51]), .C(n16919), .D(poly7_shifted[51]), .Z(n17597) );
  COND1XL U17760 ( .A(n17664), .B(n12170), .C(n17597), .Z(n10053) );
  CANR2X1 U17761 ( .A(n18028), .B(poly7_shifted[319]), .C(n17598), .D(
        poly7_shifted[307]), .Z(n17599) );
  COND1XL U17762 ( .A(n17664), .B(n18028), .C(n17599), .Z(n9797) );
  CANR2X1 U17763 ( .A(n12299), .B(poly1_shifted[62]), .C(n17714), .D(
        poly1_shifted[51]), .Z(n17600) );
  COND1XL U17764 ( .A(n17658), .B(n12299), .C(n17600), .Z(n9306) );
  CANR2X1 U17765 ( .A(n12008), .B(poly14_shifted[163]), .C(n17755), .D(
        poly14_shifted[147]), .Z(n17601) );
  COND1XL U17766 ( .A(n17664), .B(n12008), .C(n17601), .Z(n10258) );
  CIVX2 U17767 ( .A(n18176), .Z(n17654) );
  CANR2X1 U17768 ( .A(n17603), .B(poly13_shifted[353]), .C(n17613), .D(
        poly13_shifted[339]), .Z(n17602) );
  COND1XL U17769 ( .A(n17654), .B(n17603), .C(n17602), .Z(n10721) );
  CANR2X1 U17770 ( .A(n17990), .B(poly13_shifted[481]), .C(n17668), .D(
        poly13_shifted[467]), .Z(n17604) );
  COND1XL U17771 ( .A(n17654), .B(n17990), .C(n17604), .Z(n10593) );
  CANR2X1 U17772 ( .A(n17982), .B(poly13_shifted[385]), .C(poly13_shifted[371]), .D(n18017), .Z(n17605) );
  COND1XL U17773 ( .A(n17658), .B(n17982), .C(n17605), .Z(n10689) );
  CANR2X1 U17774 ( .A(n12009), .B(poly14_shifted[131]), .C(n16540), .D(
        poly14_shifted[115]), .Z(n17606) );
  COND1XL U17775 ( .A(n17664), .B(n12009), .C(n17606), .Z(n10290) );
  CANR2XL U17776 ( .A(n13124), .B(poly13_shifted[33]), .C(n17607), .D(
        poly13_shifted[19]), .Z(n17608) );
  COND1XL U17777 ( .A(n17658), .B(n13124), .C(n17608), .Z(n11041) );
  CANR2X1 U17778 ( .A(n17610), .B(poly1_shifted[158]), .C(n17458), .D(
        poly1_shifted[147]), .Z(n17609) );
  COND1XL U17779 ( .A(n17658), .B(n17610), .C(n17609), .Z(n9210) );
  CANR2X1 U17780 ( .A(n12012), .B(poly1_shifted[94]), .C(n17613), .D(
        poly1_shifted[83]), .Z(n17611) );
  COND1XL U17781 ( .A(n17658), .B(n12012), .C(n17611), .Z(n9274) );
  CANR2X1 U17782 ( .A(n13351), .B(poly9_shifted[62]), .C(n17705), .D(
        poly9_shifted[51]), .Z(n17612) );
  COND1XL U17783 ( .A(n17661), .B(n13351), .C(n17612), .Z(n11254) );
  CANR2X1 U17784 ( .A(n17615), .B(poly13_shifted[321]), .C(n17613), .D(
        poly13_shifted[307]), .Z(n17614) );
  COND1XL U17785 ( .A(n17654), .B(n17615), .C(n17614), .Z(n10753) );
  CANR2XL U17786 ( .A(n12958), .B(poly14_shifted[99]), .C(poly14_shifted[83]), 
        .D(n18017), .Z(n17616) );
  COND1XL U17787 ( .A(n17664), .B(n12958), .C(n17616), .Z(n10322) );
  CANR2X1 U17788 ( .A(n18002), .B(poly14_shifted[35]), .C(n17401), .D(
        poly14_shifted[19]), .Z(n17617) );
  COND1XL U17789 ( .A(n17658), .B(n18002), .C(n17617), .Z(n10386) );
  CANR2X1 U17790 ( .A(n16694), .B(poly14_shifted[259]), .C(n17714), .D(
        poly14_shifted[243]), .Z(n17618) );
  COND1XL U17791 ( .A(n17664), .B(n16694), .C(n17618), .Z(n10162) );
  CEOXL U17792 ( .A(Poly8[84]), .B(Poly8[69]), .Z(n17619) );
  CANR2X1 U17793 ( .A(n17750), .B(Poly8[83]), .C(n17620), .D(n17619), .Z(
        n17621) );
  COND1XL U17794 ( .A(n17661), .B(n17750), .C(n17621), .Z(n11318) );
  CANR2X1 U17795 ( .A(n17987), .B(poly13_shifted[449]), .C(n17504), .D(
        poly13_shifted[435]), .Z(n17622) );
  COND1XL U17796 ( .A(n17658), .B(n17987), .C(n17622), .Z(n10625) );
  CEOXL U17797 ( .A(Poly14[287]), .B(Poly14[195]), .Z(n17623) );
  CANR2X1 U17798 ( .A(n12202), .B(Poly14[211]), .C(n16427), .D(n17623), .Z(
        n17624) );
  COND1XL U17799 ( .A(n17664), .B(n12202), .C(n17624), .Z(n10194) );
  CEOXL U17800 ( .A(Poly12[124]), .B(Poly12[35]), .Z(n17625) );
  CANR2X1 U17801 ( .A(n12598), .B(Poly12[51]), .C(n17094), .D(n17625), .Z(
        n17626) );
  COND1XL U17802 ( .A(n17658), .B(n12598), .C(n17626), .Z(n10481) );
  CANR2X1 U17803 ( .A(n16425), .B(poly1_shifted[126]), .C(n17488), .D(
        poly1_shifted[115]), .Z(n17627) );
  COND1XL U17804 ( .A(n17658), .B(n16425), .C(n17627), .Z(n9242) );
  CENX1 U17805 ( .A(Poly11[36]), .B(n17628), .Z(n17629) );
  CANR2X1 U17806 ( .A(n17683), .B(Poly11[51]), .C(n17629), .D(n17755), .Z(
        n17630) );
  COND1XL U17807 ( .A(n17664), .B(n17683), .C(n17630), .Z(n11138) );
  CANR2X1 U17808 ( .A(n17955), .B(poly9_shifted[94]), .C(n17280), .D(
        poly9_shifted[83]), .Z(n17631) );
  COND1XL U17809 ( .A(n17661), .B(n17955), .C(n17631), .Z(n11222) );
  CANR2X1 U17810 ( .A(n18018), .B(Poly7[19]), .C(n16372), .D(poly7_shifted[19]), .Z(n17632) );
  COND1XL U17811 ( .A(n17664), .B(n18018), .C(n17632), .Z(n10085) );
  CANR2XL U17812 ( .A(n18191), .B(poly1_shifted[286]), .C(n17215), .D(
        poly1_shifted[275]), .Z(n17633) );
  COND1XL U17813 ( .A(n17658), .B(n18191), .C(n17633), .Z(n9082) );
  CANR2X1 U17814 ( .A(n17969), .B(poly13_shifted[97]), .C(n17634), .D(
        poly13_shifted[83]), .Z(n17635) );
  COND1XL U17815 ( .A(n17654), .B(n17969), .C(n17635), .Z(n10977) );
  CEOXL U17816 ( .A(Poly12[126]), .B(Poly12[67]), .Z(n17636) );
  CANR2X1 U17817 ( .A(n12161), .B(Poly12[83]), .C(n17642), .D(n17636), .Z(
        n17637) );
  COND1XL U17818 ( .A(n17658), .B(n12161), .C(n17637), .Z(n10449) );
  CENX1 U17819 ( .A(Poly8[84]), .B(Poly8[86]), .Z(n17638) );
  CENX1 U17820 ( .A(Poly8[5]), .B(n17638), .Z(n17639) );
  CANR2X1 U17821 ( .A(n12175), .B(poly8_shifted[33]), .C(n17640), .D(n17639), 
        .Z(n17641) );
  COND1XL U17822 ( .A(n17661), .B(n12175), .C(n17641), .Z(n11382) );
  CANR2X1 U17823 ( .A(n17977), .B(poly13_shifted[161]), .C(n17642), .D(
        poly13_shifted[147]), .Z(n17643) );
  COND1XL U17824 ( .A(n17658), .B(n17977), .C(n17643), .Z(n10913) );
  CANR2X1 U17825 ( .A(n17974), .B(poly13_shifted[129]), .C(n17508), .D(
        poly13_shifted[115]), .Z(n17644) );
  COND1XL U17826 ( .A(n17654), .B(n17974), .C(n17644), .Z(n10945) );
  CEOXL U17827 ( .A(Poly13[524]), .B(Poly13[165]), .Z(n17645) );
  CANR2X1 U17828 ( .A(n13014), .B(poly13_shifted[193]), .C(n16427), .D(n17645), 
        .Z(n17646) );
  COND1XL U17829 ( .A(n17658), .B(n13014), .C(n17646), .Z(n10881) );
  CANR2X1 U17830 ( .A(n12185), .B(Poly11[19]), .C(n17295), .D(
        poly11_shifted[19]), .Z(n17647) );
  COND1XL U17831 ( .A(n17664), .B(n12185), .C(n17647), .Z(n11170) );
  CANR2X1 U17832 ( .A(n12625), .B(poly7_shifted[287]), .C(n17280), .D(
        poly7_shifted[275]), .Z(n17648) );
  COND1XL U17833 ( .A(n17658), .B(n12625), .C(n17648), .Z(n9829) );
  CAN2XL U17834 ( .A(n18017), .B(poly8_shifted[51]), .Z(n17649) );
  CANR1XL U17835 ( .A(poly8_shifted[65]), .B(n12287), .C(n17649), .Z(n17650)
         );
  COND1XL U17836 ( .A(n17661), .B(n12287), .C(n17650), .Z(n11350) );
  CANR2X1 U17837 ( .A(n17652), .B(Poly12[115]), .C(n17705), .D(
        poly12_shifted[115]), .Z(n17651) );
  COND1XL U17838 ( .A(n17664), .B(n17652), .C(n17651), .Z(n10417) );
  CANR2X1 U17839 ( .A(n17491), .B(poly13_shifted[513]), .C(n17705), .D(
        poly13_shifted[499]), .Z(n17653) );
  COND1XL U17840 ( .A(n17654), .B(n17491), .C(n17653), .Z(n10561) );
  CANR2X1 U17841 ( .A(n12997), .B(Poly12[19]), .C(n17655), .D(
        poly12_shifted[19]), .Z(n17656) );
  COND1XL U17842 ( .A(n17658), .B(n12997), .C(n17656), .Z(n10513) );
  CANR2X1 U17843 ( .A(n12211), .B(Poly2[19]), .C(n17209), .D(poly2_shifted[19]), .Z(n17657) );
  COND1XL U17844 ( .A(n17658), .B(n12211), .C(n17657), .Z(n8991) );
  CANR2X1 U17845 ( .A(n12977), .B(Poly7[179]), .C(n17504), .D(
        poly7_shifted[179]), .Z(n17659) );
  COND1XL U17846 ( .A(n17664), .B(n12977), .C(n17659), .Z(n9925) );
  CANR2X1 U17847 ( .A(n17731), .B(Poly9[19]), .C(n16427), .D(poly9_shifted[19]), .Z(n17660) );
  COND1XL U17848 ( .A(n17661), .B(n17731), .C(n17660), .Z(n11286) );
  CANR2X1 U17849 ( .A(n13040), .B(poly7_shifted[351]), .C(n17285), .D(
        poly7_shifted[339]), .Z(n17662) );
  COND1XL U17850 ( .A(n17661), .B(n13040), .C(n17662), .Z(n9765) );
  CANR2X1 U17851 ( .A(n17471), .B(poly7_shifted[95]), .C(n17238), .D(
        poly7_shifted[83]), .Z(n17663) );
  COND1XL U17852 ( .A(n17664), .B(n17471), .C(n17663), .Z(n10021) );
  CANR2X1 U17853 ( .A(n12262), .B(Poly9[115]), .C(n16702), .D(
        poly9_shifted[115]), .Z(n17665) );
  COND1XL U17854 ( .A(n17658), .B(n12262), .C(n17665), .Z(n11190) );
  CANR2X1 U17855 ( .A(n17667), .B(poly13_shifted[225]), .C(n16919), .D(
        poly13_shifted[211]), .Z(n17666) );
  COND1XL U17856 ( .A(n17664), .B(n17667), .C(n17666), .Z(n10849) );
  CANR2X1 U17857 ( .A(n12900), .B(poly13_shifted[65]), .C(n17668), .D(
        poly13_shifted[51]), .Z(n17669) );
  COND1XL U17858 ( .A(n17664), .B(n12900), .C(n17669), .Z(n11009) );
  CANR2X1 U17859 ( .A(n12206), .B(poly7_shifted[383]), .C(n17094), .D(
        poly7_shifted[371]), .Z(n17670) );
  COND1XL U17860 ( .A(n17658), .B(n12206), .C(n17670), .Z(n9733) );
  CANR2X1 U17861 ( .A(n17655), .B(poly0_shifted[147]), .C(n17671), .D(
        poly0_shifted[165]), .Z(n17672) );
  COND1XL U17862 ( .A(n17674), .B(n17673), .C(n17672), .Z(n9430) );
  CENX1 U17863 ( .A(n17675), .B(Poly11[35]), .Z(n17676) );
  CANR2X1 U17864 ( .A(n17683), .B(Poly11[50]), .C(n16787), .D(n17676), .Z(
        n17677) );
  COND1XL U17865 ( .A(n17569), .B(n17683), .C(n17677), .Z(n11139) );
  CANR2X1 U17866 ( .A(n17731), .B(Poly9[18]), .C(n17705), .D(poly9_shifted[18]), .Z(n17678) );
  COND1XL U17867 ( .A(n17551), .B(n17731), .C(n17678), .Z(n11287) );
  CANR2X1 U17868 ( .A(n12262), .B(Poly9[114]), .C(n17998), .D(
        poly9_shifted[114]), .Z(n17679) );
  COND1XL U17869 ( .A(n17549), .B(n12262), .C(n17679), .Z(n11191) );
  CEOXL U17870 ( .A(n17680), .B(Poly11[19]), .Z(n17681) );
  CNR2XL U17871 ( .A(n17829), .B(n17681), .Z(n17682) );
  CANR1XL U17872 ( .A(Poly11[34]), .B(n17683), .C(n17682), .Z(n17684) );
  COND1XL U17873 ( .A(n16775), .B(n17747), .C(n17684), .Z(n11155) );
  CEOXL U17874 ( .A(Poly2[55]), .B(n17685), .Z(n17686) );
  CENX1 U17875 ( .A(Poly2[67]), .B(n17686), .Z(n17687) );
  CANR2XL U17876 ( .A(n17696), .B(Poly2[67]), .C(n17136), .D(n17687), .Z(
        n17688) );
  COND1XL U17877 ( .A(n13275), .B(n17696), .C(n17688), .Z(n8943) );
  CEOXL U17878 ( .A(Poly2[52]), .B(n17738), .Z(n17689) );
  CENX1 U17879 ( .A(Poly2[64]), .B(n17689), .Z(n17690) );
  CANR2X1 U17880 ( .A(n17696), .B(Poly2[64]), .C(n16307), .D(n17690), .Z(
        n17691) );
  COND1XL U17881 ( .A(n17751), .B(n17696), .C(n17691), .Z(n8946) );
  CEOXL U17882 ( .A(Poly2[53]), .B(n17692), .Z(n17693) );
  CENX1 U17883 ( .A(Poly2[65]), .B(n17693), .Z(n17694) );
  CANR2X1 U17884 ( .A(n17696), .B(Poly2[65]), .C(n16540), .D(n17694), .Z(
        n17695) );
  COND1XL U17885 ( .A(n17697), .B(n17696), .C(n17695), .Z(n8945) );
  CANR2X1 U17886 ( .A(n12287), .B(poly8_shifted[60]), .C(n17449), .D(
        poly8_shifted[46]), .Z(n17698) );
  COND1XL U17887 ( .A(n17699), .B(n12287), .C(n17698), .Z(n11355) );
  CENX1 U17888 ( .A(Poly8[85]), .B(Poly8[87]), .Z(n17700) );
  CENX1 U17889 ( .A(Poly8[6]), .B(n17700), .Z(n17701) );
  CANR2X1 U17890 ( .A(n12175), .B(poly8_shifted[34]), .C(n17458), .D(n17701), 
        .Z(n17702) );
  COND1XL U17891 ( .A(n17707), .B(n12175), .C(n17702), .Z(n11381) );
  CEOXL U17892 ( .A(Poly8[85]), .B(Poly8[70]), .Z(n17703) );
  CANR2XL U17893 ( .A(n17750), .B(Poly8[84]), .C(n17288), .D(n17703), .Z(
        n17704) );
  COND1XL U17894 ( .A(n17707), .B(n17750), .C(n17704), .Z(n11317) );
  CANR2X1 U17895 ( .A(n12287), .B(poly8_shifted[66]), .C(n17705), .D(
        poly8_shifted[52]), .Z(n17706) );
  COND1XL U17896 ( .A(n17707), .B(n12287), .C(n17706), .Z(n11349) );
  CANR2X1 U17897 ( .A(n12287), .B(poly8_shifted[47]), .C(n17105), .D(
        poly8_shifted[33]), .Z(n17708) );
  COND1XL U17898 ( .A(n17711), .B(n12287), .C(n17708), .Z(n11368) );
  CANR2X1 U17899 ( .A(n17955), .B(poly9_shifted[76]), .C(n17362), .D(
        poly9_shifted[65]), .Z(n17709) );
  COND1XL U17900 ( .A(n17711), .B(n17955), .C(n17709), .Z(n11240) );
  CANR2X1 U17901 ( .A(n17731), .B(poly9_shifted[12]), .C(n17375), .D(
        Poly9[106]), .Z(n17710) );
  COND1XL U17902 ( .A(n17711), .B(n17731), .C(n17710), .Z(n11304) );
  CEOXL U17903 ( .A(Poly9[113]), .B(Poly9[92]), .Z(n17712) );
  CANR2X1 U17904 ( .A(n12262), .B(poly9_shifted[114]), .C(n17755), .D(n17712), 
        .Z(n17713) );
  COND1XL U17905 ( .A(n17718), .B(n12262), .C(n17713), .Z(n11202) );
  CANR2X1 U17906 ( .A(n12175), .B(Poly8[7]), .C(n17714), .D(Poly8[89]), .Z(
        n17715) );
  COND1XL U17907 ( .A(n17718), .B(n12175), .C(n17715), .Z(n11394) );
  CANR2X1 U17908 ( .A(n13351), .B(poly9_shifted[50]), .C(n16583), .D(
        poly9_shifted[39]), .Z(n17716) );
  COND1XL U17909 ( .A(n17718), .B(n13351), .C(n17716), .Z(n11266) );
  CANR2X1 U17910 ( .A(n17955), .B(poly9_shifted[82]), .C(n18234), .D(
        poly9_shifted[71]), .Z(n17717) );
  COND1XL U17911 ( .A(n17718), .B(n17955), .C(n17717), .Z(n11234) );
  CANR2X1 U17912 ( .A(n12287), .B(poly8_shifted[70]), .C(n17174), .D(
        poly8_shifted[56]), .Z(n17719) );
  COND1XL U17913 ( .A(n17721), .B(n12287), .C(n17719), .Z(n11345) );
  CANR2X1 U17914 ( .A(n17955), .B(Poly9[88]), .C(n17158), .D(poly9_shifted[88]), .Z(n17720) );
  COND1XL U17915 ( .A(n17721), .B(n17955), .C(n17720), .Z(n11217) );
  CANR2X1 U17916 ( .A(n12287), .B(poly8_shifted[69]), .C(n17755), .D(
        poly8_shifted[55]), .Z(n17722) );
  COND1XL U17917 ( .A(n12296), .B(n12287), .C(n17722), .Z(n11346) );
  CANR2X1 U17918 ( .A(n17955), .B(Poly9[87]), .C(n17343), .D(poly9_shifted[87]), .Z(n17723) );
  COND1XL U17919 ( .A(n12000), .B(n17955), .C(n17723), .Z(n11218) );
  CANR2X1 U17920 ( .A(n13351), .B(poly9_shifted[66]), .C(n17755), .D(
        poly9_shifted[55]), .Z(n17724) );
  COND1XL U17921 ( .A(n12296), .B(n13351), .C(n17724), .Z(n11250) );
  CANR2X1 U17922 ( .A(n12185), .B(Poly11[23]), .C(n16479), .D(
        poly11_shifted[23]), .Z(n17725) );
  COND1XL U17923 ( .A(n12000), .B(n12185), .C(n17725), .Z(n11166) );
  CANR2X1 U17924 ( .A(n12185), .B(Poly11[28]), .C(n17174), .D(
        poly11_shifted[28]), .Z(n17726) );
  COND1XL U17925 ( .A(n11978), .B(n12185), .C(n17726), .Z(n11161) );
  CANR2X1 U17926 ( .A(n12185), .B(poly11_shifted[24]), .C(n17209), .D(
        Poly11[80]), .Z(n17727) );
  COND1XL U17927 ( .A(n12002), .B(n12185), .C(n17727), .Z(n11180) );
  CANR2X1 U17928 ( .A(n12287), .B(poly8_shifted[55]), .C(n17755), .D(
        poly8_shifted[41]), .Z(n17728) );
  COND1XL U17929 ( .A(n12002), .B(n12287), .C(n17728), .Z(n11360) );
  CANR2XL U17930 ( .A(n17731), .B(poly9_shifted[20]), .C(Poly9[114]), .D(
        n18017), .Z(n17729) );
  COND1XL U17931 ( .A(n12002), .B(n17731), .C(n17729), .Z(n11296) );
  CANR2X1 U17932 ( .A(n17731), .B(poly9_shifted[16]), .C(n17215), .D(
        Poly9[110]), .Z(n17730) );
  COND1XL U17933 ( .A(n11981), .B(n17731), .C(n17730), .Z(n11300) );
  CANR2X1 U17934 ( .A(n17955), .B(Poly9[90]), .C(n17280), .D(poly9_shifted[90]), .Z(n17733) );
  COND1XL U17935 ( .A(n17735), .B(n17955), .C(n17733), .Z(n11215) );
  CANR2X1 U17936 ( .A(n12161), .B(Poly12[90]), .C(n17998), .D(
        poly12_shifted[90]), .Z(n17734) );
  COND1XL U17937 ( .A(n17735), .B(n12161), .C(n17734), .Z(n10442) );
  CANR2X1 U17938 ( .A(n12185), .B(Poly11[26]), .C(n17390), .D(
        poly11_shifted[26]), .Z(n17736) );
  COND1XL U17939 ( .A(n17735), .B(n12185), .C(n17736), .Z(n11163) );
  CANR2X1 U17940 ( .A(n17750), .B(Poly8[72]), .C(n17504), .D(poly8_shifted[72]), .Z(n17737) );
  COND1XL U17941 ( .A(n17163), .B(n17750), .C(n17737), .Z(n11329) );
  CENX1 U17942 ( .A(Poly2[47]), .B(n17738), .Z(n17739) );
  CANR2X1 U17943 ( .A(n17306), .B(Poly2[59]), .C(n17458), .D(n17739), .Z(
        n17740) );
  COND1XL U17944 ( .A(n17741), .B(n17306), .C(n17740), .Z(n8951) );
  CEOXL U17945 ( .A(Poly11[17]), .B(n17742), .Z(n17743) );
  CNR2XL U17946 ( .A(n17744), .B(n17743), .Z(n17745) );
  CANR1XL U17947 ( .A(Poly11[32]), .B(n17747), .C(n17745), .Z(n17746) );
  COND1XL U17948 ( .A(n17751), .B(n17747), .C(n17746), .Z(n11157) );
  CANR2X1 U17949 ( .A(n17935), .B(poly5_shifted[46]), .C(n17545), .D(
        poly5_shifted[32]), .Z(n17748) );
  COND1XL U17950 ( .A(n17751), .B(n17935), .C(n17748), .Z(n11494) );
  CANR2X1 U17951 ( .A(n17750), .B(poly8_shifted[78]), .C(n17466), .D(
        poly8_shifted[64]), .Z(n17749) );
  COND1XL U17952 ( .A(n17751), .B(n17750), .C(n17749), .Z(n11337) );
  CANR2X1 U17953 ( .A(n13351), .B(poly9_shifted[65]), .C(n17755), .D(
        poly9_shifted[54]), .Z(n17752) );
  COND1XL U17954 ( .A(n17753), .B(n13351), .C(n17752), .Z(n11251) );
  CANR2X1 U17955 ( .A(n13351), .B(poly9_shifted[49]), .C(n16307), .D(
        poly9_shifted[38]), .Z(n17754) );
  COND1XL U17956 ( .A(n17757), .B(n13351), .C(n17754), .Z(n11267) );
  CANR2X1 U17957 ( .A(n12175), .B(Poly8[6]), .C(n17755), .D(Poly8[88]), .Z(
        n17756) );
  COND1XL U17958 ( .A(n17757), .B(n12175), .C(n17756), .Z(n11395) );
  CNR2IXL U17959 ( .B(datain[5]), .A(n17799), .Z(n17758) );
  CANR1X1 U17960 ( .A(entrophy[5]), .B(n17759), .C(n17758), .Z(n17762) );
  CAN3X1 U17961 ( .A(n17762), .B(n17761), .C(n17760), .Z(n17764) );
  CANR11X1 U17962 ( .A(n17766), .B(n17765), .C(n17764), .D(n17763), .Z(n17819)
         );
  CND2XL U17963 ( .A(n17768), .B(n17767), .Z(n17772) );
  CANR1XL U17964 ( .A(n17770), .B(datain[6]), .C(n17769), .Z(n17771) );
  CANR11X1 U17965 ( .A(n17773), .B(n17772), .C(n17771), .D(n14977), .Z(n17818)
         );
  CAOR2X1 U17966 ( .A(n17775), .B(entrophy[22]), .C(entrophy[26]), .D(n17774), 
        .Z(n17783) );
  CND2XL U17967 ( .A(n17776), .B(entrophy[15]), .Z(n17781) );
  CIVXL U17968 ( .A(n17777), .Z(n17780) );
  CANR11X1 U17969 ( .A(n17781), .B(n17780), .C(n17779), .D(n17778), .Z(n17782)
         );
  CNR2X1 U17970 ( .A(n17783), .B(n17782), .Z(n17789) );
  CNR3XL U17971 ( .A(n17785), .B(n14226), .C(n17784), .Z(n17786) );
  CANR1XL U17972 ( .A(n17787), .B(entrophy[17]), .C(n17786), .Z(n17788) );
  CND2X1 U17973 ( .A(n17789), .B(n17788), .Z(n17817) );
  CIVXL U17974 ( .A(n17790), .Z(n17796) );
  CANR1XL U17975 ( .A(datain[7]), .B(n17792), .C(n17791), .Z(n17795) );
  CAN4X1 U17976 ( .A(n17796), .B(n17795), .C(n17794), .D(n17793), .Z(n17815)
         );
  CNR2X1 U17977 ( .A(n17797), .B(entrophy[12]), .Z(n17803) );
  CNR2XL U17978 ( .A(entrophy[7]), .B(dataselector[47]), .Z(n17798) );
  CANR4CX1 U17979 ( .A(n17803), .B(n17802), .C(n17801), .D(n17800), .Z(n17811)
         );
  COND1XL U17980 ( .A(entrophy[21]), .B(n17805), .C(n17804), .Z(n17806) );
  CANR3X1 U17981 ( .A(n17809), .B(n17808), .C(n17807), .D(n17806), .Z(n17810)
         );
  CANR3X1 U17982 ( .A(scrambler[15]), .B(n17959), .C(n17811), .D(n17810), .Z(
        n17814) );
  CANR2X1 U17983 ( .A(n17812), .B(entrophy[18]), .C(entrophy[11]), .D(n11971), 
        .Z(n17813) );
  COND3X1 U17984 ( .A(n17815), .B(n12055), .C(n17814), .D(n17813), .Z(n17816)
         );
  COR4X1 U17985 ( .A(n17819), .B(n17818), .C(n17817), .D(n17816), .Z(n8715) );
  CENX1 U17986 ( .A(dataselector[2]), .B(n17821), .Z(n17822) );
  CENX1 U17987 ( .A(n17822), .B(dataselector[61]), .Z(n17827) );
  CIVX1 U17988 ( .A(dataselector[9]), .Z(n17823) );
  CNR2XL U17989 ( .A(n17831), .B(n17823), .Z(n17824) );
  CANR1XL U17990 ( .A(n18189), .B(n17832), .C(n17824), .Z(n17825) );
  COND1XL U17991 ( .A(n17827), .B(n17826), .C(n17825), .Z(n8786) );
  CENX1 U17992 ( .A(polydata[1]), .B(scrambler[24]), .Z(n17833) );
  CENX1 U17993 ( .A(n17834), .B(n17833), .Z(dataout[14]) );
  CEOXL U17994 ( .A(scrambler[19]), .B(n17921), .Z(n17836) );
  CENX1 U17995 ( .A(polydata[3]), .B(scrambler[26]), .Z(n17835) );
  CENX1 U17996 ( .A(n17836), .B(n17835), .Z(dataout[12]) );
  CENX1 U17997 ( .A(scrambler[9]), .B(scrambler[21]), .Z(n17837) );
  CENX1 U17998 ( .A(n17838), .B(n17837), .Z(n17840) );
  CENX1 U17999 ( .A(scrambler[23]), .B(n17891), .Z(n17839) );
  CENX1 U18000 ( .A(n17840), .B(n17839), .Z(dataout[25]) );
  CEOX1 U18001 ( .A(scrambler[23]), .B(scrambler[25]), .Z(n17899) );
  CENX1 U18002 ( .A(scrambler[27]), .B(n17899), .Z(n17886) );
  CENX1 U18003 ( .A(polydata[9]), .B(n17912), .Z(n17841) );
  CENX1 U18004 ( .A(n17842), .B(n17841), .Z(n17843) );
  CEOX1 U18005 ( .A(n17880), .B(n17843), .Z(n17844) );
  CENX1 U18006 ( .A(n17886), .B(n17844), .Z(dataout[6]) );
  CEOX1 U18007 ( .A(n17921), .B(n17911), .Z(n17846) );
  CENX1 U18008 ( .A(scrambler[2]), .B(scrambler[29]), .Z(n17845) );
  CENX1 U18009 ( .A(n17846), .B(n17845), .Z(dataout[18]) );
  CEOX1 U18010 ( .A(scrambler[19]), .B(scrambler[20]), .Z(n17888) );
  CEOX1 U18011 ( .A(n17888), .B(n17871), .Z(n17848) );
  CENX1 U18012 ( .A(scrambler[11]), .B(scrambler[17]), .Z(n17847) );
  CENX1 U18013 ( .A(n17848), .B(n17847), .Z(dataout[27]) );
  CENX1 U18014 ( .A(n17888), .B(scrambler[18]), .Z(n17849) );
  CENX1 U18015 ( .A(n17886), .B(n17849), .Z(n17850) );
  CENX1 U18016 ( .A(polydata[2]), .B(n17850), .Z(dataout[13]) );
  CEOX1 U18017 ( .A(n17868), .B(n17851), .Z(n17853) );
  CEOX1 U18018 ( .A(n17880), .B(n17899), .Z(n17895) );
  CENX1 U18019 ( .A(polydata[15]), .B(n17895), .Z(n17852) );
  CENX1 U18020 ( .A(n17853), .B(n17852), .Z(dataout[0]) );
  CEOX1 U18021 ( .A(n17899), .B(n17854), .Z(n17857) );
  CEOX1 U18022 ( .A(scrambler[21]), .B(n17857), .Z(n17856) );
  CENX1 U18023 ( .A(polydata[4]), .B(scrambler[31]), .Z(n17855) );
  CENX1 U18024 ( .A(n17856), .B(n17855), .Z(dataout[11]) );
  CEOX1 U18025 ( .A(n17857), .B(n17907), .Z(n17859) );
  CENX1 U18026 ( .A(scrambler[0]), .B(scrambler[24]), .Z(n17858) );
  CENX1 U18027 ( .A(n17859), .B(n17858), .Z(dataout[16]) );
  CEOXL U18028 ( .A(scrambler[26]), .B(scrambler[23]), .Z(n17876) );
  CEOX1 U18029 ( .A(n17876), .B(n17893), .Z(n17861) );
  CENX1 U18030 ( .A(n17907), .B(scrambler[8]), .Z(n17860) );
  CENX1 U18031 ( .A(n17861), .B(n17860), .Z(dataout[24]) );
  CENX1 U18032 ( .A(n17907), .B(n17891), .Z(n17865) );
  CEOX1 U18033 ( .A(n17862), .B(n17865), .Z(n17864) );
  CENX1 U18034 ( .A(scrambler[6]), .B(scrambler[18]), .Z(n17863) );
  CENX1 U18035 ( .A(n17864), .B(n17863), .Z(dataout[22]) );
  CEOX1 U18036 ( .A(n17865), .B(n17868), .Z(n17867) );
  CENX1 U18037 ( .A(polydata[5]), .B(scrambler[28]), .Z(n17866) );
  CENX1 U18038 ( .A(n17867), .B(n17866), .Z(dataout[10]) );
  CENX1 U18039 ( .A(n17868), .B(n17905), .Z(n17869) );
  CENX1 U18040 ( .A(n17883), .B(n17869), .Z(n17870) );
  CENX1 U18041 ( .A(polydata[0]), .B(n17870), .Z(dataout[15]) );
  CEOX1 U18042 ( .A(scrambler[7]), .B(n17871), .Z(n17873) );
  CENX1 U18043 ( .A(scrambler[31]), .B(scrambler[22]), .Z(n17872) );
  CENX1 U18044 ( .A(n17873), .B(n17872), .Z(n17874) );
  CENX1 U18045 ( .A(n17874), .B(n17883), .Z(dataout[23]) );
  CEOXL U18046 ( .A(n17876), .B(n17875), .Z(n17878) );
  CENX1 U18047 ( .A(n17884), .B(scrambler[5]), .Z(n17877) );
  CENX1 U18048 ( .A(n17878), .B(n17877), .Z(n17879) );
  CEOX1 U18049 ( .A(n17880), .B(n17879), .Z(n17881) );
  CENX1 U18050 ( .A(n17882), .B(n17881), .Z(dataout[21]) );
  CENX1 U18051 ( .A(n17884), .B(n17883), .Z(n17910) );
  CENX1 U18052 ( .A(scrambler[31]), .B(n17910), .Z(n17885) );
  CENX1 U18053 ( .A(n17886), .B(n17885), .Z(n17887) );
  CENX1 U18054 ( .A(polydata[7]), .B(n17887), .Z(dataout[8]) );
  CENX1 U18055 ( .A(n17889), .B(n17888), .Z(n17890) );
  CENX1 U18056 ( .A(n17891), .B(n17890), .Z(n17892) );
  CENX1 U18057 ( .A(polydata[8]), .B(n17892), .Z(dataout[7]) );
  CENX1 U18058 ( .A(n17893), .B(n17912), .Z(n17896) );
  CENX1 U18059 ( .A(scrambler[3]), .B(scrambler[30]), .Z(n17894) );
  CENX1 U18060 ( .A(n17896), .B(n17894), .Z(dataout[19]) );
  CEOX1 U18061 ( .A(n17896), .B(n17895), .Z(n17898) );
  CENX1 U18062 ( .A(n17907), .B(scrambler[12]), .Z(n17897) );
  CENX1 U18063 ( .A(n17898), .B(n17897), .Z(dataout[28]) );
  CEOX1 U18064 ( .A(scrambler[31]), .B(scrambler[17]), .Z(n17902) );
  CEOX1 U18065 ( .A(n17902), .B(n17899), .Z(n17901) );
  CENX1 U18066 ( .A(polydata[10]), .B(scrambler[26]), .Z(n17900) );
  CENX1 U18067 ( .A(n17901), .B(n17900), .Z(dataout[5]) );
  CENX1 U18068 ( .A(n17902), .B(n17912), .Z(n17906) );
  CENX1 U18069 ( .A(scrambler[28]), .B(scrambler[21]), .Z(n17920) );
  CENX1 U18070 ( .A(scrambler[27]), .B(n17920), .Z(n17923) );
  CEOX1 U18071 ( .A(n17906), .B(n17923), .Z(n17904) );
  CENX1 U18072 ( .A(polydata[13]), .B(scrambler[22]), .Z(n17903) );
  CENX1 U18073 ( .A(n17904), .B(n17903), .Z(dataout[2]) );
  CEOX1 U18074 ( .A(n17906), .B(n17905), .Z(n17909) );
  CENX1 U18075 ( .A(n17907), .B(scrambler[14]), .Z(n17908) );
  CENX1 U18076 ( .A(n17909), .B(n17908), .Z(dataout[30]) );
  CEOX1 U18077 ( .A(n17911), .B(n17910), .Z(n17914) );
  CENX1 U18078 ( .A(scrambler[24]), .B(n17912), .Z(n17918) );
  CENX1 U18079 ( .A(scrambler[13]), .B(n17918), .Z(n17913) );
  CENX1 U18080 ( .A(n17914), .B(n17913), .Z(dataout[29]) );
  CEOXL U18081 ( .A(scrambler[1]), .B(scrambler[17]), .Z(n17916) );
  CENX1 U18082 ( .A(scrambler[29]), .B(scrambler[23]), .Z(n17915) );
  CENX1 U18083 ( .A(n17916), .B(n17915), .Z(n17917) );
  CEOX1 U18084 ( .A(n17918), .B(n17917), .Z(n17919) );
  CENX1 U18085 ( .A(n17920), .B(n17919), .Z(dataout[17]) );
  CENX1 U18086 ( .A(scrambler[15]), .B(n17921), .Z(n17922) );
  CENX1 U18087 ( .A(n17923), .B(n17922), .Z(dataout[31]) );
  CANR1XL U18088 ( .A(n17925), .B(n17924), .C(n16381), .Z(n17929) );
  CANR2X1 U18089 ( .A(n17930), .B(poly5_shifted[25]), .C(n17926), .D(
        Poly5[122]), .Z(n17927) );
  COND1XL U18090 ( .A(n17929), .B(n17928), .C(n17927), .Z(n11515) );
  COND1XL U18091 ( .A(poly5_shifted[25]), .B(n17934), .C(n18196), .Z(n17933)
         );
  CND2X1 U18092 ( .A(n17930), .B(poly5_shifted[39]), .Z(n17931) );
  COND1XL U18093 ( .A(n17933), .B(n17932), .C(n17931), .Z(n11501) );
  COND1XL U18094 ( .A(poly5_shifted[57]), .B(n17934), .C(n18196), .Z(n17937)
         );
  CND2X1 U18095 ( .A(n17935), .B(poly5_shifted[71]), .Z(n17936) );
  COND1XL U18096 ( .A(n17937), .B(n15378), .C(n17936), .Z(n11469) );
  CANR1XL U18097 ( .A(n17939), .B(n17938), .C(n12007), .Z(n17943) );
  CANR2XL U18098 ( .A(n17942), .B(Poly5[92]), .C(n17940), .D(Poly5[78]), .Z(
        n17941) );
  COND1XL U18099 ( .A(n17943), .B(n17942), .C(n17941), .Z(n11434) );
  COND1XL U18100 ( .A(poly8_shifted[34]), .B(n12415), .C(n18126), .Z(n17945)
         );
  CND2X1 U18101 ( .A(n12287), .B(poly8_shifted[48]), .Z(n17944) );
  COND1XL U18102 ( .A(n17945), .B(n12287), .C(n17944), .Z(n11367) );
  COND1XL U18103 ( .A(poly8_shifted[37]), .B(n11994), .C(n18134), .Z(n17947)
         );
  CND2X1 U18104 ( .A(n12287), .B(poly8_shifted[51]), .Z(n17946) );
  COND1XL U18105 ( .A(n17947), .B(n12287), .C(n17946), .Z(n11364) );
  COND1XL U18106 ( .A(poly8_shifted[47]), .B(n18206), .C(n18163), .Z(n17949)
         );
  CND2X1 U18107 ( .A(n12287), .B(poly8_shifted[61]), .Z(n17948) );
  COND1XL U18108 ( .A(n17949), .B(n12287), .C(n17948), .Z(n11354) );
  COND1XL U18109 ( .A(poly8_shifted[50]), .B(n18210), .C(n18172), .Z(n17951)
         );
  CND2X1 U18110 ( .A(n12287), .B(poly8_shifted[64]), .Z(n17950) );
  COND1XL U18111 ( .A(n17951), .B(n12287), .C(n17950), .Z(n11351) );
  COND1XL U18112 ( .A(poly9_shifted[67]), .B(n18053), .C(n18111), .Z(n17953)
         );
  CND2X1 U18113 ( .A(n17955), .B(poly9_shifted[78]), .Z(n17952) );
  COND1XL U18114 ( .A(n17953), .B(n17955), .C(n17952), .Z(n11238) );
  COND1XL U18115 ( .A(poly9_shifted[79]), .B(n18206), .C(n18163), .Z(n17956)
         );
  CND2X1 U18116 ( .A(n17955), .B(poly9_shifted[90]), .Z(n17954) );
  COND1XL U18117 ( .A(n17956), .B(n17955), .C(n17954), .Z(n11226) );
  CIVX1 U18118 ( .A(Poly10[3]), .Z(n17958) );
  CANR1XL U18119 ( .A(n17957), .B(n17958), .C(n18206), .Z(n17963) );
  CNR3XL U18120 ( .A(n17959), .B(Poly10[41]), .C(n17958), .Z(n17960) );
  CANR1XL U18121 ( .A(Poly10[15]), .B(n17962), .C(n17960), .Z(n17961) );
  COND1XL U18122 ( .A(n17963), .B(n17962), .C(n17961), .Z(n11088) );
  CND2X1 U18123 ( .A(n12003), .B(n17964), .Z(n18183) );
  CANR2X1 U18124 ( .A(n17965), .B(poly13_shifted[63]), .C(poly13_shifted[77]), 
        .D(n12900), .Z(n17966) );
  COND1XL U18125 ( .A(n17967), .B(n18183), .C(n17966), .Z(n10997) );
  COND1XL U18126 ( .A(poly13_shifted[86]), .B(n18034), .C(n18088), .Z(n17970)
         );
  CND2X1 U18127 ( .A(n17969), .B(poly13_shifted[100]), .Z(n17968) );
  COND1XL U18128 ( .A(n17970), .B(n17969), .C(n17968), .Z(n10974) );
  COND1XL U18129 ( .A(poly13_shifted[110]), .B(n18160), .C(n18159), .Z(n17972)
         );
  CND2X1 U18130 ( .A(n17974), .B(poly13_shifted[124]), .Z(n17971) );
  COND1XL U18131 ( .A(n17972), .B(n17974), .C(n17971), .Z(n10950) );
  COND1XL U18132 ( .A(poly13_shifted[127]), .B(n12003), .C(n18022), .Z(n17975)
         );
  CND2X1 U18133 ( .A(n17974), .B(poly13_shifted[141]), .Z(n17973) );
  COND1XL U18134 ( .A(n17975), .B(n17974), .C(n17973), .Z(n10933) );
  COND1XL U18135 ( .A(poly13_shifted[154]), .B(n18095), .C(n18094), .Z(n17978)
         );
  CND2X1 U18136 ( .A(n17977), .B(poly13_shifted[168]), .Z(n17976) );
  COND1XL U18137 ( .A(n17978), .B(n17977), .C(n17976), .Z(n10906) );
  COND1XL U18138 ( .A(poly13_shifted[352]), .B(n12010), .C(n18185), .Z(n17980)
         );
  CND2X1 U18139 ( .A(n17982), .B(poly13_shifted[366]), .Z(n17979) );
  COND1XL U18140 ( .A(n17980), .B(n17982), .C(n17979), .Z(n10708) );
  COND1XL U18141 ( .A(poly13_shifted[365]), .B(n18219), .C(n18156), .Z(n17983)
         );
  CND2X1 U18142 ( .A(n17982), .B(poly13_shifted[379]), .Z(n17981) );
  COND1XL U18143 ( .A(n17983), .B(n17982), .C(n17981), .Z(n10695) );
  COND1XL U18144 ( .A(poly13_shifted[425]), .B(n18189), .C(n18188), .Z(n17985)
         );
  CND2X1 U18145 ( .A(n17987), .B(poly13_shifted[439]), .Z(n17984) );
  COND1XL U18146 ( .A(n17985), .B(n17987), .C(n17984), .Z(n10635) );
  COND1XL U18147 ( .A(poly13_shifted[432]), .B(n18167), .C(n18166), .Z(n17988)
         );
  CND2X1 U18148 ( .A(n17987), .B(poly13_shifted[446]), .Z(n17986) );
  COND1XL U18149 ( .A(n17988), .B(n17987), .C(n17986), .Z(n10628) );
  COND1XL U18150 ( .A(poly13_shifted[450]), .B(n12415), .C(n18126), .Z(n17991)
         );
  CND2X1 U18151 ( .A(n17990), .B(poly13_shifted[464]), .Z(n17989) );
  COND1XL U18152 ( .A(n17991), .B(n17990), .C(n17989), .Z(n10610) );
  COND1XL U18153 ( .A(poly12_shifted[24]), .B(n13994), .C(n18091), .Z(n17993)
         );
  CND2X1 U18154 ( .A(n12997), .B(Poly12[24]), .Z(n17992) );
  COND1XL U18155 ( .A(n17993), .B(n12997), .C(n17992), .Z(n10508) );
  COND1XL U18156 ( .A(poly12_shifted[62]), .B(n18105), .C(n18104), .Z(n17997)
         );
  CND2X1 U18157 ( .A(n12598), .B(Poly12[62]), .Z(n17996) );
  COND1XL U18158 ( .A(n17997), .B(n12598), .C(n17996), .Z(n10470) );
  CANR2XL U18159 ( .A(n18001), .B(n11999), .C(n17998), .D(poly12_shifted[119]), 
        .Z(n17999) );
  COND1XL U18160 ( .A(n18001), .B(n18000), .C(n17999), .Z(n10413) );
  CANR2X1 U18161 ( .A(n17280), .B(poly14_shifted[31]), .C(poly14_shifted[47]), 
        .D(n18002), .Z(n18003) );
  COND1XL U18162 ( .A(n18004), .B(n18183), .C(n18003), .Z(n10374) );
  COND1XL U18163 ( .A(poly14_shifted[73]), .B(n18189), .C(n18188), .Z(n18006)
         );
  CND2X1 U18164 ( .A(n12958), .B(poly14_shifted[89]), .Z(n18005) );
  COND1XL U18165 ( .A(n18006), .B(n12958), .C(n18005), .Z(n10332) );
  COND1XL U18166 ( .A(poly14_shifted[78]), .B(n18160), .C(n18159), .Z(n18008)
         );
  CND2X1 U18167 ( .A(n12958), .B(poly14_shifted[94]), .Z(n18007) );
  COND1XL U18168 ( .A(n18008), .B(n12958), .C(n18007), .Z(n10327) );
  COND1XL U18169 ( .A(poly14_shifted[200]), .B(n18142), .C(n18141), .Z(n18010)
         );
  CND2X1 U18170 ( .A(n12202), .B(Poly14[200]), .Z(n18009) );
  COND1XL U18171 ( .A(n18010), .B(n12202), .C(n18009), .Z(n10205) );
  COND1XL U18172 ( .A(poly14_shifted[234]), .B(n12013), .C(n18147), .Z(n18012)
         );
  CND2X1 U18173 ( .A(n16694), .B(poly14_shifted[250]), .Z(n18011) );
  COND1XL U18174 ( .A(n18012), .B(n16694), .C(n18011), .Z(n10171) );
  COND1XL U18175 ( .A(poly14_shifted[242]), .B(n18210), .C(n18172), .Z(n18014)
         );
  CND2X1 U18176 ( .A(n16694), .B(poly14_shifted[258]), .Z(n18013) );
  COND1XL U18177 ( .A(n18014), .B(n16694), .C(n18013), .Z(n10163) );
  COND1XL U18178 ( .A(poly14_shifted[264]), .B(n18142), .C(n18141), .Z(n18016)
         );
  CND2X1 U18179 ( .A(n12932), .B(poly14_shifted[280]), .Z(n18015) );
  COND1XL U18180 ( .A(n18016), .B(n12932), .C(n18015), .Z(n10141) );
  COND1XL U18181 ( .A(poly7_shifted[158]), .B(n18105), .C(n18104), .Z(n18021)
         );
  CND2X1 U18182 ( .A(n13070), .B(poly7_shifted[170]), .Z(n18020) );
  COND1XL U18183 ( .A(n18021), .B(n13070), .C(n18020), .Z(n9946) );
  COND1XL U18184 ( .A(poly7_shifted[159]), .B(n14436), .C(n18022), .Z(n18024)
         );
  CND2X1 U18185 ( .A(n13070), .B(poly7_shifted[171]), .Z(n18023) );
  COND1XL U18186 ( .A(n18024), .B(n13070), .C(n18023), .Z(n9945) );
  COND1XL U18187 ( .A(poly7_shifted[164]), .B(n12004), .C(n18131), .Z(n18026)
         );
  CND2X1 U18188 ( .A(n12977), .B(poly7_shifted[176]), .Z(n18025) );
  COND1XL U18189 ( .A(n18026), .B(n12977), .C(n18025), .Z(n9940) );
  COND1XL U18190 ( .A(poly7_shifted[290]), .B(n12415), .C(n18126), .Z(n18029)
         );
  CND2X1 U18191 ( .A(n18028), .B(poly7_shifted[302]), .Z(n18027) );
  COND1XL U18192 ( .A(n18029), .B(n18028), .C(n18027), .Z(n9814) );
  COND1XL U18193 ( .A(poly7_shifted[330]), .B(n12013), .C(n18147), .Z(n18031)
         );
  CND2X1 U18194 ( .A(n13040), .B(poly7_shifted[342]), .Z(n18030) );
  COND1XL U18195 ( .A(n18031), .B(n13040), .C(n18030), .Z(n9774) );
  COND1XL U18196 ( .A(Poly15[47]), .B(n12415), .C(n18126), .Z(n18033) );
  CND2X1 U18197 ( .A(n18044), .B(poly15_shifted[17]), .Z(n18032) );
  COND1XL U18198 ( .A(n18033), .B(n18044), .C(n18032), .Z(n9635) );
  COND1XL U18199 ( .A(poly15_shifted[22]), .B(n18034), .C(n18088), .Z(n18036)
         );
  CND2X1 U18200 ( .A(n18044), .B(Poly15[22]), .Z(n18035) );
  COND1XL U18201 ( .A(n18036), .B(n18044), .C(n18035), .Z(n9615) );
  COND1XL U18202 ( .A(poly15_shifted[25]), .B(n18249), .C(n18196), .Z(n18038)
         );
  CND2X1 U18203 ( .A(n18044), .B(Poly15[25]), .Z(n18037) );
  COND1XL U18204 ( .A(n18038), .B(n18044), .C(n18037), .Z(n9612) );
  CEOX1 U18205 ( .A(Poly15[13]), .B(Poly15[45]), .Z(n18041) );
  COAN1XL U18206 ( .A(n18040), .B(n18041), .C(n11978), .Z(n18045) );
  CANR2X1 U18207 ( .A(n18044), .B(Poly15[28]), .C(n18042), .D(n18041), .Z(
        n18043) );
  COND1XL U18208 ( .A(n18045), .B(n18044), .C(n18043), .Z(n9609) );
  CANR2X1 U18209 ( .A(n16565), .B(n18048), .C(n18047), .D(poly15_shifted[49]), 
        .Z(n18049) );
  COND1XL U18210 ( .A(n16565), .B(n18050), .C(n18049), .Z(n9588) );
  COND1XL U18211 ( .A(poly0_shifted[64]), .B(n12010), .C(n18185), .Z(n18052)
         );
  CND2X1 U18212 ( .A(n12291), .B(poly0_shifted[82]), .Z(n18051) );
  COND1XL U18213 ( .A(n18052), .B(n12291), .C(n18051), .Z(n9513) );
  COND1XL U18214 ( .A(poly0_shifted[67]), .B(n18053), .C(n18111), .Z(n18055)
         );
  CND2X1 U18215 ( .A(n12291), .B(poly0_shifted[85]), .Z(n18054) );
  COND1XL U18216 ( .A(n18055), .B(n12291), .C(n18054), .Z(n9510) );
  COND1XL U18217 ( .A(poly0_shifted[68]), .B(n12004), .C(n18131), .Z(n18057)
         );
  CND2X1 U18218 ( .A(n12291), .B(poly0_shifted[86]), .Z(n18056) );
  COND1XL U18219 ( .A(n18057), .B(n12291), .C(n18056), .Z(n9509) );
  COND1XL U18220 ( .A(poly0_shifted[72]), .B(n18142), .C(n18141), .Z(n18059)
         );
  CND2X1 U18221 ( .A(n12291), .B(poly0_shifted[90]), .Z(n18058) );
  COND1XL U18222 ( .A(n18059), .B(n12291), .C(n18058), .Z(n9505) );
  COND1XL U18223 ( .A(poly0_shifted[73]), .B(n18189), .C(n18188), .Z(n18061)
         );
  CND2X1 U18224 ( .A(n12291), .B(poly0_shifted[91]), .Z(n18060) );
  COND1XL U18225 ( .A(n18061), .B(n12291), .C(n18060), .Z(n9504) );
  COND1XL U18226 ( .A(poly0_shifted[74]), .B(n12013), .C(n18147), .Z(n18063)
         );
  CND2X1 U18227 ( .A(n12291), .B(poly0_shifted[92]), .Z(n18062) );
  COND1XL U18228 ( .A(n18063), .B(n12291), .C(n18062), .Z(n9503) );
  COND1XL U18229 ( .A(poly0_shifted[75]), .B(n16381), .C(n18150), .Z(n18065)
         );
  CND2X1 U18230 ( .A(n12291), .B(poly0_shifted[93]), .Z(n18064) );
  COND1XL U18231 ( .A(n18065), .B(n12291), .C(n18064), .Z(n9502) );
  COND1XL U18232 ( .A(poly0_shifted[76]), .B(n13028), .C(n18153), .Z(n18067)
         );
  CND2X1 U18233 ( .A(n12291), .B(poly0_shifted[94]), .Z(n18066) );
  COND1XL U18234 ( .A(n18067), .B(n12291), .C(n18066), .Z(n9501) );
  COND1XL U18235 ( .A(poly0_shifted[77]), .B(n18219), .C(n18156), .Z(n18069)
         );
  CND2X1 U18236 ( .A(n12291), .B(poly0_shifted[95]), .Z(n18068) );
  COND1XL U18237 ( .A(n18069), .B(n12291), .C(n18068), .Z(n9500) );
  COND1XL U18238 ( .A(poly0_shifted[78]), .B(n18160), .C(n18159), .Z(n18071)
         );
  CND2X1 U18239 ( .A(n12291), .B(poly0_shifted[96]), .Z(n18070) );
  COND1XL U18240 ( .A(n18071), .B(n12291), .C(n18070), .Z(n9499) );
  COND1XL U18241 ( .A(poly0_shifted[79]), .B(n18206), .C(n18163), .Z(n18073)
         );
  CND2X1 U18242 ( .A(n12291), .B(poly0_shifted[97]), .Z(n18072) );
  COND1XL U18243 ( .A(n18073), .B(n12291), .C(n18072), .Z(n9498) );
  COND1XL U18244 ( .A(poly0_shifted[80]), .B(n12381), .C(n18166), .Z(n18075)
         );
  CND2X1 U18245 ( .A(n12291), .B(poly0_shifted[98]), .Z(n18074) );
  COND1XL U18246 ( .A(n18075), .B(n12291), .C(n18074), .Z(n9497) );
  COND1XL U18247 ( .A(n13522), .B(poly0_shifted[81]), .C(n18193), .Z(n18077)
         );
  CND2X1 U18248 ( .A(n12291), .B(poly0_shifted[99]), .Z(n18076) );
  COND1XL U18249 ( .A(n18077), .B(n12291), .C(n18076), .Z(n9496) );
  COND1XL U18250 ( .A(poly0_shifted[82]), .B(n18210), .C(n18172), .Z(n18079)
         );
  CND2X1 U18251 ( .A(n12291), .B(poly0_shifted[100]), .Z(n18078) );
  COND1XL U18252 ( .A(n18079), .B(n12291), .C(n18078), .Z(n9495) );
  COND1XL U18253 ( .A(poly0_shifted[83]), .B(n18176), .C(n18175), .Z(n18081)
         );
  CND2X1 U18254 ( .A(n12291), .B(poly0_shifted[101]), .Z(n18080) );
  COND1XL U18255 ( .A(n18081), .B(n12291), .C(n18080), .Z(n9494) );
  COND1XL U18256 ( .A(poly0_shifted[84]), .B(n18082), .C(n18200), .Z(n18084)
         );
  CND2X1 U18257 ( .A(n12291), .B(poly0_shifted[102]), .Z(n18083) );
  COND1XL U18258 ( .A(n18084), .B(n12291), .C(n18083), .Z(n9493) );
  COND1XL U18259 ( .A(poly0_shifted[85]), .B(n18241), .C(n18085), .Z(n18087)
         );
  CND2X1 U18260 ( .A(n12291), .B(poly0_shifted[103]), .Z(n18086) );
  COND1XL U18261 ( .A(n18087), .B(n12291), .C(n18086), .Z(n9492) );
  COND1XL U18262 ( .A(poly0_shifted[86]), .B(n14487), .C(n18088), .Z(n18090)
         );
  CND2X1 U18263 ( .A(n12291), .B(poly0_shifted[104]), .Z(n18089) );
  COND1XL U18264 ( .A(n18090), .B(n12291), .C(n18089), .Z(n9491) );
  COND1XL U18265 ( .A(poly0_shifted[88]), .B(n13994), .C(n18091), .Z(n18093)
         );
  CND2X1 U18266 ( .A(n12291), .B(poly0_shifted[106]), .Z(n18092) );
  COND1XL U18267 ( .A(n18093), .B(n12291), .C(n18092), .Z(n9489) );
  COND1XL U18268 ( .A(poly0_shifted[90]), .B(n18095), .C(n18094), .Z(n18097)
         );
  CND2X1 U18269 ( .A(n12291), .B(poly0_shifted[108]), .Z(n18096) );
  COND1XL U18270 ( .A(n18097), .B(n12291), .C(n18096), .Z(n9487) );
  COND1XL U18271 ( .A(poly0_shifted[91]), .B(n18099), .C(n18098), .Z(n18101)
         );
  CND2X1 U18272 ( .A(n12291), .B(poly0_shifted[109]), .Z(n18100) );
  COND1XL U18273 ( .A(n18101), .B(n12291), .C(n18100), .Z(n9486) );
  COND1XL U18274 ( .A(poly0_shifted[92]), .B(n12007), .C(n18224), .Z(n18103)
         );
  CND2X1 U18275 ( .A(n12291), .B(poly0_shifted[110]), .Z(n18102) );
  COND1XL U18276 ( .A(n18103), .B(n12291), .C(n18102), .Z(n9485) );
  COND1XL U18277 ( .A(poly0_shifted[94]), .B(n18105), .C(n18104), .Z(n18107)
         );
  CND2X1 U18278 ( .A(n12291), .B(poly0_shifted[112]), .Z(n18106) );
  COND1XL U18279 ( .A(n18107), .B(n12291), .C(n18106), .Z(n9483) );
  COND1XL U18280 ( .A(poly0_shifted[192]), .B(n18108), .C(n18185), .Z(n18110)
         );
  CND2XL U18281 ( .A(n18119), .B(poly0_shifted[210]), .Z(n18109) );
  COND1XL U18282 ( .A(n18110), .B(n18119), .C(n18109), .Z(n9385) );
  COND1XL U18283 ( .A(poly0_shifted[195]), .B(n18053), .C(n18111), .Z(n18113)
         );
  CND2XL U18284 ( .A(n18119), .B(poly0_shifted[213]), .Z(n18112) );
  COND1XL U18285 ( .A(n18113), .B(n18119), .C(n18112), .Z(n9382) );
  COND1XL U18286 ( .A(poly0_shifted[196]), .B(n12004), .C(n18131), .Z(n18115)
         );
  CND2XL U18287 ( .A(n18119), .B(poly0_shifted[214]), .Z(n18114) );
  COND1XL U18288 ( .A(n18115), .B(n18119), .C(n18114), .Z(n9381) );
  COND1XL U18289 ( .A(poly0_shifted[201]), .B(n18189), .C(n18188), .Z(n18120)
         );
  CND2XL U18290 ( .A(n18119), .B(poly0_shifted[219]), .Z(n18118) );
  COND1XL U18291 ( .A(n18120), .B(n18119), .C(n18118), .Z(n9376) );
  COND1XL U18292 ( .A(Poly1[336]), .B(n12010), .C(n18185), .Z(n18122) );
  CND2XL U18293 ( .A(n18180), .B(poly1_shifted[11]), .Z(n18121) );
  COND1XL U18294 ( .A(n18122), .B(n18180), .C(n18121), .Z(n9357) );
  COND1XL U18295 ( .A(Poly1[337]), .B(n12020), .C(n18123), .Z(n18125) );
  CND2XL U18296 ( .A(n18180), .B(poly1_shifted[12]), .Z(n18124) );
  COND1XL U18297 ( .A(n18125), .B(n18180), .C(n18124), .Z(n9356) );
  COND1XL U18298 ( .A(Poly1[338]), .B(n12415), .C(n18126), .Z(n18128) );
  CND2XL U18299 ( .A(n18180), .B(poly1_shifted[13]), .Z(n18127) );
  COND1XL U18300 ( .A(n18128), .B(n18180), .C(n18127), .Z(n9355) );
  CND2XL U18301 ( .A(n18180), .B(poly1_shifted[14]), .Z(n18129) );
  COND1XL U18302 ( .A(n18130), .B(n18180), .C(n18129), .Z(n9354) );
  COND1XL U18303 ( .A(Poly1[340]), .B(n12004), .C(n18131), .Z(n18133) );
  CND2XL U18304 ( .A(n18180), .B(poly1_shifted[15]), .Z(n18132) );
  COND1XL U18305 ( .A(n18133), .B(n18180), .C(n18132), .Z(n9353) );
  COND1XL U18306 ( .A(Poly1[341]), .B(n11984), .C(n18134), .Z(n18136) );
  CND2XL U18307 ( .A(n18180), .B(poly1_shifted[16]), .Z(n18135) );
  COND1XL U18308 ( .A(n18136), .B(n18180), .C(n18135), .Z(n9352) );
  COND1XL U18309 ( .A(Poly1[343]), .B(n18138), .C(n18137), .Z(n18140) );
  CND2XL U18310 ( .A(n18180), .B(poly1_shifted[18]), .Z(n18139) );
  COND1XL U18311 ( .A(n18140), .B(n18180), .C(n18139), .Z(n9350) );
  COND1XL U18312 ( .A(Poly1[344]), .B(n18142), .C(n18141), .Z(n18144) );
  CND2XL U18313 ( .A(n18180), .B(poly1_shifted[19]), .Z(n18143) );
  COND1XL U18314 ( .A(n18144), .B(n18180), .C(n18143), .Z(n9349) );
  COND1XL U18315 ( .A(Poly1[345]), .B(n18189), .C(n18188), .Z(n18146) );
  CND2XL U18316 ( .A(n18180), .B(poly1_shifted[20]), .Z(n18145) );
  COND1XL U18317 ( .A(n18146), .B(n18180), .C(n18145), .Z(n9348) );
  COND1XL U18318 ( .A(Poly1[346]), .B(n12013), .C(n18147), .Z(n18149) );
  CND2XL U18319 ( .A(n18180), .B(poly1_shifted[21]), .Z(n18148) );
  COND1XL U18320 ( .A(n18149), .B(n18180), .C(n18148), .Z(n9347) );
  COND1XL U18321 ( .A(poly1_shifted[11]), .B(n16381), .C(n18150), .Z(n18152)
         );
  CND2XL U18322 ( .A(n18180), .B(poly1_shifted[22]), .Z(n18151) );
  COND1XL U18323 ( .A(n18152), .B(n18180), .C(n18151), .Z(n9346) );
  COND1XL U18324 ( .A(poly1_shifted[12]), .B(n13028), .C(n18153), .Z(n18155)
         );
  CND2XL U18325 ( .A(n18180), .B(poly1_shifted[23]), .Z(n18154) );
  COND1XL U18326 ( .A(n18155), .B(n18180), .C(n18154), .Z(n9345) );
  COND1XL U18327 ( .A(poly1_shifted[13]), .B(n18219), .C(n18156), .Z(n18158)
         );
  CND2XL U18328 ( .A(n18180), .B(poly1_shifted[24]), .Z(n18157) );
  COND1XL U18329 ( .A(n18158), .B(n18180), .C(n18157), .Z(n9344) );
  COND1XL U18330 ( .A(poly1_shifted[14]), .B(n18160), .C(n18159), .Z(n18162)
         );
  CND2XL U18331 ( .A(n18180), .B(poly1_shifted[25]), .Z(n18161) );
  COND1XL U18332 ( .A(n18162), .B(n18180), .C(n18161), .Z(n9343) );
  COND1XL U18333 ( .A(poly1_shifted[15]), .B(n18206), .C(n18163), .Z(n18165)
         );
  CND2XL U18334 ( .A(n18180), .B(poly1_shifted[26]), .Z(n18164) );
  COND1XL U18335 ( .A(n18165), .B(n18180), .C(n18164), .Z(n9342) );
  COND1XL U18336 ( .A(poly1_shifted[16]), .B(n18167), .C(n18166), .Z(n18169)
         );
  CND2XL U18337 ( .A(n18180), .B(poly1_shifted[27]), .Z(n18168) );
  COND1XL U18338 ( .A(n18169), .B(n18180), .C(n18168), .Z(n9341) );
  COND1XL U18339 ( .A(n18048), .B(poly1_shifted[17]), .C(n18193), .Z(n18171)
         );
  CND2XL U18340 ( .A(n18180), .B(poly1_shifted[28]), .Z(n18170) );
  COND1XL U18341 ( .A(n18171), .B(n18180), .C(n18170), .Z(n9340) );
  COND1XL U18342 ( .A(poly1_shifted[18]), .B(n18210), .C(n18172), .Z(n18174)
         );
  CND2XL U18343 ( .A(n18180), .B(poly1_shifted[29]), .Z(n18173) );
  COND1XL U18344 ( .A(n18174), .B(n18180), .C(n18173), .Z(n9339) );
  COND1XL U18345 ( .A(poly1_shifted[19]), .B(n18176), .C(n18175), .Z(n18178)
         );
  CND2XL U18346 ( .A(n18180), .B(poly1_shifted[30]), .Z(n18177) );
  COND1XL U18347 ( .A(n18178), .B(n18180), .C(n18177), .Z(n9338) );
  CENX1 U18348 ( .A(Poly1[336]), .B(n18179), .Z(n18181) );
  CANR2XL U18349 ( .A(n17280), .B(n18181), .C(poly1_shifted[42]), .D(n18180), 
        .Z(n18182) );
  COND1XL U18350 ( .A(n18184), .B(n18183), .C(n18182), .Z(n9326) );
  COND1XL U18351 ( .A(poly1_shifted[96]), .B(n12010), .C(n18185), .Z(n18187)
         );
  CND2X1 U18352 ( .A(n16425), .B(poly1_shifted[107]), .Z(n18186) );
  COND1XL U18353 ( .A(n18187), .B(n16425), .C(n18186), .Z(n9261) );
  COND1XL U18354 ( .A(poly1_shifted[265]), .B(n18189), .C(n18188), .Z(n18192)
         );
  CND2X1 U18355 ( .A(n18191), .B(poly1_shifted[276]), .Z(n18190) );
  COND1XL U18356 ( .A(n18192), .B(n18191), .C(n18190), .Z(n9092) );
  COND1XL U18357 ( .A(n13522), .B(poly1_shifted[305]), .C(n18193), .Z(n18195)
         );
  CND2X1 U18358 ( .A(n18198), .B(poly1_shifted[316]), .Z(n18194) );
  COND1XL U18359 ( .A(n18195), .B(n18198), .C(n18194), .Z(n9052) );
  COND1XL U18360 ( .A(poly1_shifted[313]), .B(n18249), .C(n18196), .Z(n18199)
         );
  CND2X1 U18361 ( .A(n18198), .B(poly1_shifted[324]), .Z(n18197) );
  COND1XL U18362 ( .A(n18199), .B(n18198), .C(n18197), .Z(n9044) );
  COND1XL U18363 ( .A(poly3_shifted[20]), .B(n18082), .C(n18200), .Z(n18202)
         );
  CND2X1 U18364 ( .A(n15737), .B(poly3_shifted[34]), .Z(n18201) );
  COND1XL U18365 ( .A(n18202), .B(n15737), .C(n18201), .Z(n8920) );
  COND1XL U18366 ( .A(poly3_shifted[23]), .B(n11999), .C(n18203), .Z(n18205)
         );
  CND2X1 U18367 ( .A(n15737), .B(poly3_shifted[37]), .Z(n18204) );
  COND1XL U18368 ( .A(n18205), .B(n15737), .C(n18204), .Z(n8917) );
  CANR2X1 U18369 ( .A(n18206), .B(n18209), .C(n16985), .D(poly3_shifted[79]), 
        .Z(n18207) );
  COND1XL U18370 ( .A(n18208), .B(n18212), .C(n18207), .Z(n8861) );
  CANR2XL U18371 ( .A(n18210), .B(n18209), .C(n17285), .D(poly3_shifted[82]), 
        .Z(n18211) );
  COND1XL U18372 ( .A(n18213), .B(n18212), .C(n18211), .Z(n8858) );
  CANR1XL U18373 ( .A(n18214), .B(n18220), .C(n16381), .Z(n18217) );
  CIVXL U18374 ( .A(n18214), .Z(n18215) );
  CANR2X1 U18375 ( .A(n18230), .B(poly4_shifted[28]), .C(n18221), .D(n18215), 
        .Z(n18216) );
  COND1XL U18376 ( .A(n18217), .B(n18230), .C(n18216), .Z(n8845) );
  COND1XL U18377 ( .A(n18220), .B(n18219), .C(n18218), .Z(n18223) );
  CANR2X1 U18378 ( .A(n18230), .B(poly4_shifted[30]), .C(n18221), .D(Poly4[59]), .Z(n18222) );
  COND1XL U18379 ( .A(n18230), .B(n18223), .C(n18222), .Z(n8843) );
  COND1XL U18380 ( .A(poly4_shifted[28]), .B(n12007), .C(n18224), .Z(n18226)
         );
  CND2X1 U18381 ( .A(n18230), .B(Poly4[28]), .Z(n18225) );
  COND1XL U18382 ( .A(n18226), .B(n18230), .C(n18225), .Z(n8828) );
  COND1XL U18383 ( .A(poly4_shifted[29]), .B(n18228), .C(n18227), .Z(n18231)
         );
  CND2X1 U18384 ( .A(n18230), .B(Poly4[29]), .Z(n18229) );
  COND1XL U18385 ( .A(n18231), .B(n18230), .C(n18229), .Z(n8827) );
  CEOXL U18386 ( .A(dataselector[62]), .B(dataselector[27]), .Z(n18232) );
  CENX1 U18387 ( .A(n18233), .B(n18232), .Z(n18235) );
  CANR2X1 U18388 ( .A(n18235), .B(n18234), .C(n12415), .D(n18248), .Z(n18236)
         );
  COND1XL U18389 ( .A(n18252), .B(n18237), .C(n18236), .Z(n8761) );
  CENX1 U18390 ( .A(n18239), .B(n18238), .Z(n18240) );
  CENX1 U18391 ( .A(dataselector[46]), .B(n18240), .Z(n18242) );
  CANR2X1 U18392 ( .A(n18242), .B(n17508), .C(n18241), .D(n18248), .Z(n18243)
         );
  COND1XL U18393 ( .A(n18244), .B(n18252), .C(n18243), .Z(n8742) );
  CENX1 U18394 ( .A(n18245), .B(dataselector[50]), .Z(n18246) );
  CENX1 U18395 ( .A(n18247), .B(n18246), .Z(n18250) );
  CANR2X1 U18396 ( .A(n18250), .B(n17094), .C(n18249), .D(n18248), .Z(n18251)
         );
  COND1XL U18397 ( .A(n18253), .B(n18252), .C(n18251), .Z(n8738) );
endmodule

