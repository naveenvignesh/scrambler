`timescale 1ns/10ps
module scrambler_serialin_mux(clk,rst,pd_sel,p0,p1,p2,p3,p4,p5,p6,p7,p8,p9,p10,p11,p12,p13,p14,p15,polydataout);

input             clk,rst;
input  [4:0]       pd_sel;        
input  [220-1:0]   p0;
input  [347-1:0]   p1;
input  [70 -1:0]   p2;
input  [84 -1:0]   p3;
input  [61 -1:0]   p4;
input  [125-1:0]   p5;
input  [56 -1:0]   p6;
input  [411-1:0]   p7;
input  [96 -1:0]   p8;
input  [116-1:0]   p9;
input  [43 -1:0]   p10;
input  [86 -1:0]   p11;
input  [127-1:0]   p12;
input  [528-1:0]   p13;
input  [301-1:0]   p14;
input  [60 -1:0]   p15;
output [15:0]    polydataout;


reg [15:0] polydata;


assign polydataout = rst ? 16'b0:polydata;


always@(*) begin
  
  case(pd_sel)
  0:polydata = {p0[110] ,p9[24]  ,p13[113],p14[162],p10[20],p8[17] ,p4[21]  ,p5[35] ,p1[120] ,p11[25],p2[36] ,p7[278] ,p6[15] ,p12[17] ,p15[54],p3[13]  }; 
  1:polydata = {p9[91]  ,p13[299],p10[39] ,p15[14] ,p3[42] ,p8[76] ,p7[146] ,p4[30] ,p1[116] ,p5[20] ,p6[41] ,p14[117],p0[184],p2[16]  ,p11[49],p12[90] };
  2:polydata = {p2[34]  ,p6[28]  ,p7[92]  ,p13[67] ,p9[60] ,p1[71] ,p14[52] ,p8[59] ,p4[45]  ,p15[33],p5[10] ,p3[63]  ,p10[2] ,p12[108],p11[71],p0[116] };
  3:polydata = {p14[253],p13[487],p9[69]  ,p7[178] ,p11[73],p6[33] ,p5[19]  ,p15[16],p3[25]  ,p4[14] ,p8[90] ,p10[1]  ,p12[97],p1[248] ,p0[93] ,p2[17]  }; 
  4:polydata = {p1[302] ,p4[12]  ,p13[418],p12[95] ,p5[79] ,p2[37] ,p9[38]  ,p15[35],p10[41] ,p8[36] ,p7[337],p6[53]  ,p3[69] ,p0[145] ,p11[67],p14[198]};
  5:polydata = {p9[94]  ,p0[50]  ,p14[102],p2[24]  ,p11[28],p4[19] ,p6[17]  ,p1[61] ,p12[106],p8[73] ,p7[349],p3[28]  ,p5[112],p13[338],p15[31],p10[14] };
  6:polydata = {p9[80]  ,p7[368] ,p6[21]  ,p4[25]  ,p11[72],p1[90] ,p10[11] ,p2[1]  ,p3[81]  ,p8[63] ,p15[21],p14[177],p0[52] ,p5[80]  ,p12[64],p13[219]}; 
  7:polydata = {p13[206],p3[60]  ,p9[22]  ,p5[114] ,p10[4] ,p2[43] ,p14[231],p4[38] ,p12[73] ,p0[200],p11[32],p1[249] ,p6[11] ,p15[32] ,p7[307],p8[21]  };   
  8:polydata = {p1[178] ,p6[48]  ,p12[0]  ,p8[33]  ,p7[318],p13[72],p2[26]  ,p14[62],p0[190] ,p4[57] ,p5[85] ,p15[10] ,p11[61],p9[23]  ,p10[27],p3[67]  };
  9:polydata = {p4[26] ,p11[39] ,p14[184],p8[2],p15[7],p0[173],p3[1],p12[91],p2[25],p7[73],p13[479],p6[0],p5[49],p9[33],p1[294],p10[33]     }; 
 10:polydata = {p7[222],p1[264],p12[16],p6[20],p2[30],p13[268],p9[97],p10[12] ,p14[281],p4[23],p5[38],p11[53],p0[207],p8[54],p3[53],p15[55] };  
 11:polydata = {p14[59],p1[295],p4[49],p10[10],p12[42],p11[84],p15[17],p8[52] ,p13[11],p6[43],p3[31],p7[187],p9[37],p2[38],p0[128],p5[36]   };   
 12:polydata = {p8[3],p13[351],p1[149],p14[155],p10[25],p6[54],p9[3],p15[12],p2[58],p4[37],p3[32],p11[46],p12[28],p5[43],p7[46],p0[139]     };
 13:polydata = {p13[274],p7[40],p8[67],p10[6],p0[101],p11[23],p14[248],p6[25] ,p4[11],p9[89],p12[46],p3[9],p2[4],p15[27],p1[134],p5[5]      };   
 14:polydata = {p8[64],p12[43],p5[31],p10[15],p3[57],p1[319],p6[51],p9[44],p11[81],p13[385],p15[9],p0[123],p14[192],p2[50],p4[39],p7[6]	  };     
 15:polydata = {p4[51],p2[60],p5[52],p14[61],p11[40],p8[41],p13[443],p9[65],p0[34],p15[13],p3[58],p1[300],p7[134],p12[115],p10[18],p6[24]	  };  
 16:polydata = {p7[212],p1[236],p0[156],p5[12],p2[65],p13[119],p3[71],p12[31],p11[74],p15[46],p9[68],p4[4],p10[32],p6[16],p14[226],p8[23]   };    	
 17:polydata = {p15[48],p1[244],p9[56],p5[68],p2[69],p10[37],p7[25],p6[14],p12[29],p4[32],p0[176],p3[8],p8[8],p13[411],p11[21],p14[273]     };    				
 18:polydata = {p3[7],p13[266],p9[57],p1[245],p5[122],p15[5],p7[310],p8[18],p10[31],p6[1],p2[62],p11[43],p14[237],p4[16],p12[4],p0[125]	  };   
 19:polydata = {p11[11],p3[49],p4[9],p0[178],p8[68],p5[62],p2[68],p7[320],p13[394],p1[103],p15[8],p12[68],p10[13],p6[42],p14[75],p9[40]	  };   
 20:polydata = {p13[481],p1[163],p14[194],p0[69],p11[63],p9[42],p6[8],p12[58],p7[147],p8[30],p10[38],p4[33],p2[46],p3[82],p15[58],p5[11]	  };   
 21:polydata = {p2[31],p1[70],p7[90],p12[27],p13[96],p10[28],p15[49],p5[8],p3[22],p6[29],p11[38],p14[49],p0[194],p8[44],p4[47],p9[41]	  };   
 22:polydata = {p9[93],p4[54],p6[26],p5[44],p13[493],p8[45],p15[24],p14[154],p1[222],p2[8],p12[38],p7[267],p11[14],p3[39],p10[3],p0[71]	  };   
 23:polydata = {p7[67],p6[27],p2[67],p8[22],p5[86],p15[28],p9[11],p14[139],p12[72],p4[34],p1[89],p10[34],p11[0],p13[376],p0[212],p3[3]	  };   
 24:polydata = {p14[57],p8[20],p7[378],p11[35],p5[117],p12[119],p6[7],p0[199] ,p3[41],p10[22],p9[17],p15[0],p13[436],p2[13],p4[8],p1[166]	  };   
 25:polydata = {p2[63],p3[61],p9[49],p14[218],p4[20],p15[15],p5[113],p7[152],p11[68],p1[339],p13[151],p0[109],p6[50],p10[8],p12[8],p8[24]	  };   
 26:polydata = {p6[32],p11[54],p7[140],p3[65],p15[57],p0[11],p10[7],p9[76],p5[26],p14[50],p1[307],p12[7],p13[174],p4[44],p2[54],p8[39]	  };   
 27:polydata = {p15[40],p9[101],p5[82],p11[78],p2[11],p13[506],p14[210],p0[211],p6[19],p1[304],p7[398],p4[35],p10[16],p8[61],p12[32],p3[46] };   	
 28:polydata = {p12[54],p7[218],p2[41],p6[12],p11[9],p13[241],p4[2],p9[100],p1[85],p10[5],p14[153],p3[79],p15[59],p5[24],p0[146],p8[1]	  };   
 29:polydata = {p10[0],p7[367],p12[110],p13[140],p5[74],p0[181],p4[48],p1[254],p15[47],p6[18],p11[17],p9[78],p8[25],p14[35],p2[5],p3[6]  	  };   	
 30:polydata = {p2[21],p10[30],p4[58],p3[30],p6[45],p15[37],p11[36],p9[31],p1[36],p7[47],p8[74],p12[3],p0[197],p14[285],p5[97],p13[524]	  };   
 31:polydata = {p7[118],p5[22],p1[284],p9[48],p8[58],p13[212],p3[77],p14[205] ,p6[4],p0[31],p2[44],p12[74],p4[22],p11[83],p15[45],p10[40]	  };   	
  
  endcase

end 


endmodule 

