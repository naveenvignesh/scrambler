`timescale 1ns/10ps
module scrambler_initial_load(clk,rst,datain,entrophy,scramble_sel,scramble_load);
input         clk,rst;
input  [7:0]  datain;
input  [31:0] entrophy;
input  [4:0]  scramble_sel;
output [31:0] scramble_load;

reg    [31:0] load;
assign scramble_load = rst ? 32'b0: load;


always@(*) begin 
             load =0;
      case(scramble_sel)
          0 :load =    {datain[7],entrophy[8],entrophy[1],entrophy[15],entrophy[25],entrophy[22],entrophy[7],datain[0],entrophy[19],entrophy[31],datain[3],datain[1],entrophy[29],entrophy[28],entrophy[4],datain[5],entrophy[26],entrophy[17],entrophy[11],entrophy[23],datain[2],datain[4],entrophy[13],entrophy[3],entrophy[30],entrophy[6],entrophy[9],entrophy[21],entrophy[2],entrophy[27],entrophy[18],datain[6]};
          1 :load =    {entrophy[8],entrophy[24],entrophy[7],entrophy[13],entrophy[25],entrophy[11],entrophy[21],entrophy[17],entrophy[6],entrophy[2],datain[1],entrophy[1],datain[6] ,entrophy[16],datain[0],entrophy[18],entrophy[15],entrophy[31],datain[3],datain[4],entrophy[27],entrophy[30],datain[5],entrophy[20],entrophy[28],entrophy[0],entrophy[23],datain[7],entrophy[12],entrophy[19],entrophy[14],datain[2] };
          2 :load =    {datain[4],datain[6],entrophy[2],datain[0],entrophy[24],entrophy[16],datain[7],entrophy[4],entrophy[19],entrophy[0],entrophy[28],entrophy[7] ,entrophy[20],entrophy[13],entrophy[6],datain[5],entrophy[17],entrophy[26],entrophy[30],entrophy[10],datain[1],entrophy[8],entrophy[25],entrophy[31],entrophy[22],entrophy[9],entrophy[5],entrophy[1],datain[3],entrophy[12],entrophy[3],datain[2]};
          3 :load =    {datain[1],entrophy[29],entrophy[22],datain[7],datain[4],entrophy[17],datain[2],entrophy[5],entrophy[30],datain[5],entrophy[24] ,entrophy[31],entrophy[14],entrophy[0],entrophy[6],entrophy[9],entrophy[18],datain[6],entrophy[4],entrophy[20],entrophy[27],entrophy[3],entrophy[11],entrophy[12 ],entrophy[2],entrophy[10],entrophy[25],entrophy[23],datain[0],datain[3],entrophy[21],entrophy[15]};
          4 :load =    {entrophy[6],datain[0],datain[2],entrophy[8],entrophy[29],entrophy[9],datain[5],datain[6],datain[1],entrophy[3],entrophy[14] ,entrophy[12],entrophy[17],entrophy[27],entrophy[7],entrophy[28],datain[4],datain[3],entrophy[5],entrophy[23],entrophy[0],entrophy[11],entrophy[24],entrophy[4],entrophy[1],entrophy[21],entrophy[18],entrophy[2],entrophy[22],entrophy[31],entrophy[10],datain[7]};
          5 :load =    {entrophy[18],entrophy[28],entrophy[17],entrophy[10],entrophy[14],entrophy[5],entrophy[2],datain[1],entrophy[27],entrophy[23],entrophy[31],datain[7] ,datain[0],datain[2],entrophy[21],datain[4],entrophy[7],datain[3],entrophy[11],entrophy[12],entrophy[3],entrophy[9],entrophy[15],entrophy[19],datain[6],entrophy[6],entrophy[8],entrophy[26],entrophy[0],datain[5],entrophy[29],entrophy[1]};
          6 :load =    {entrophy[30],entrophy[12],entrophy[9],entrophy[18],entrophy[16],entrophy[4],entrophy[23],entrophy[0],entrophy[1],datain[4],datain[0],datain[7] ,entrophy[27],entrophy[20],entrophy[25],entrophy[24],datain[3],datain[5],entrophy[10],entrophy[13],entrophy[6],entrophy[31],datain[2],entrophy[15],entrophy[21],entrophy[14],entrophy[26],datain[1],entrophy[3],entrophy[2],datain[6],entrophy[19]};  
          7 :load =    {datain[7],entrophy[14],entrophy[3],entrophy[24],entrophy[15],entrophy[0],entrophy[22],datain[1],entrophy[16],entrophy[8],entrophy[5],entrophy[27] ,entrophy[13],datain[3],datain[6],datain[4],datain[5],entrophy[31],datain[0],entrophy[2],entrophy[17],entrophy[4],entrophy[18],entrophy[7],entrophy[19],entrophy[1],datain[2],entrophy[6],entrophy[9],entrophy[29],entrophy[12],entrophy[25]};
          8 :load =   {datain[7],entrophy[7],entrophy[4],entrophy[1],entrophy[12],entrophy[0],entrophy[18],datain[4],datain[3],datain[5],datain[6] ,entrophy[5],entrophy[29],entrophy[17],entrophy[22],datain[0],entrophy[30],entrophy[20],entrophy[19],entrophy[13],entrophy[24],entrophy[2],datain[2],entrophy[3],entrophy[16],datain[1],entrophy[6],entrophy[15],entrophy[27],entrophy[26],entrophy[21],entrophy[23]};
          9 :load =   {entrophy[30],datain[5],entrophy[8],entrophy[20],entrophy[24],entrophy[11],entrophy[14],entrophy[1],entrophy[17],entrophy[26],entrophy[15],entrophy[16] ,datain[7],entrophy[3],entrophy[22],entrophy[13],entrophy[6],entrophy[23],entrophy[31],entrophy[7],entrophy[12],entrophy[28],datain[0],entrophy[5],datain[6],datain[4],entrophy[0],entrophy[25],datain[3],datain[1],datain[2],entrophy[18]};
         10 :load =   {entrophy[8],datain[4],entrophy[4],entrophy[6],entrophy[13],entrophy[15],entrophy[20],entrophy[10],entrophy[30],entrophy[28],datain[0],entrophy[26] ,datain[7],entrophy[16],datain[5],entrophy[19],entrophy[11],entrophy[5],entrophy[24],datain[2],entrophy[31],entrophy[25],entrophy[7],datain[1],entrophy[23],entrophy[12],datain[6],entrophy[9],entrophy[14],entrophy[21],entrophy[3],datain[3]};
         11 :load =   {entrophy[18],entrophy[27],entrophy[2],entrophy[10],entrophy[12],entrophy[28],entrophy[29],entrophy[16],datain[3],entrophy[0],entrophy[21],entrophy[26] ,datain[4],entrophy[30],datain[5],datain[1],entrophy[22],entrophy[13],datain[2],datain[7],entrophy[15],entrophy[11] ,entrophy[25],datain[0],entrophy[31],entrophy[17],datain[6],entrophy[24],entrophy[14],entrophy[23],entrophy[20],entrophy[5]};
         12 :load =   {datain[1],datain[5],entrophy[2],entrophy[5],entrophy[4],entrophy[29],entrophy[7],datain[0],entrophy[30],entrophy[26],datain[7],entrophy[15] ,entrophy[9],entrophy[27],datain[2],entrophy[25],entrophy[0],entrophy[8],entrophy[16],datain[3],entrophy[22],entrophy[6],entrophy[23],entrophy[31],entrophy[11],entrophy[19],datain[4],entrophy[24],datain[6],entrophy[17],entrophy[21],entrophy[1]};
         13 :load =   {entrophy[27],entrophy[31],entrophy[0],entrophy[1],entrophy[26],entrophy[25],entrophy[9],entrophy[23],entrophy[10],datain[0],entrophy[12],entrophy[4],entrophy[29] ,entrophy[5],entrophy[15],datain[3],entrophy[21],datain[1],entrophy[14],datain[4],entrophy[16],entrophy[3],entrophy[20],entrophy[30],entrophy[8],datain[6],entrophy[18],entrophy[2],datain[5],datain[2],datain[7],entrophy[19]};
         14 :load =   {entrophy[0],entrophy[4],entrophy[8],entrophy[3],entrophy[26],entrophy[13],entrophy[15],datain[7],entrophy[21],datain[0],entrophy[14],entrophy[28] ,datain[6],entrophy[6],entrophy[16],datain[2],entrophy[10],entrophy[1],entrophy[17],entrophy[18],entrophy[5],datain[3],entrophy[7],datain[ 4],datain[1],entrophy[29],entrophy[11],entrophy[12],entrophy[22],entrophy[2],datain[5],entrophy[19]};
         15 :load =   {datain[3],entrophy[24],datain[7],entrophy[7],datain[6],entrophy[3],entrophy[1],datain[1],entrophy[4],entrophy[11],entrophy[6],datain[0] ,entrophy[5],entrophy[23],entrophy[20],entrophy[27],datain[2],entrophy[19],entrophy[0],entrophy[26],entrophy[13],entrophy[2],entrophy[17],datain[5],entrophy[29],entrophy[8],entrophy[31],entrophy[18],entrophy[16],datain[4],entrophy[21],entrophy[9]};
         16 :load =   {entrophy[30],entrophy[22],entrophy[26],entrophy[17],entrophy[31],entrophy[25],entrophy[8],datain[4],entrophy[14],entrophy[10],entrophy[29],datain[5] ,entrophy[18],entrophy[27],entrophy[13],datain[6],datain[2],entrophy[9],entrophy[16],entrophy[20],datain[1],entrophy[24],entrophy[15],entrophy[4],datain[0],entrophy[19],entrophy[2],datain[7],entrophy[5],entrophy[1],datain[3],entrophy[7]};
         17 :load =   {entrophy[21],entrophy[8],entrophy[11],entrophy[9],datain[2],entrophy[16],datain[4],entrophy[1],datain[0],entrophy[30],entrophy[13],entrophy[27] ,entrophy[20],datain[7],entrophy[23],datain[3],datain[6],entrophy[12],entrophy[19],entrophy[15],entrophy[14],entrophy[29],entrophy[0],datain[1],entrophy[24],entrophy[5],entrophy[22],entrophy[3],entrophy[2],entrophy[28],entrophy[7],datain[5]};
         18 :load =    {entrophy[0],entrophy[27],entrophy[20],entrophy[3],entrophy[29],entrophy[22],datain[5],entrophy[8],datain[4],entrophy[4],entrophy[11],entrophy[31] ,datain[7],entrophy[2],entrophy[7],entrophy[9],datain[2],datain[6],datain[0],datain[3],entrophy[1],entrophy[25],entrophy[19],datain[1],entrophy[13],entrophy[21],entrophy[28],entrophy[30],entrophy[18],entrophy[14],entrophy[26],entrophy[24] };
         19 :load =   {entrophy[10],entrophy[28],entrophy[30],entrophy[3],datain[2],entrophy[22],entrophy[29],datain[5],entrophy[0],entrophy[16],entrophy[17],entrophy[6] ,entrophy[15],datain[6],entrophy[8],entrophy[1],entrophy[5],entrophy[4],entrophy[9],entrophy[2],entrophy[27],entrophy[13],datain[1],entrophy[7],entrophy[18 ],datain[4],datain[0],datain[3],entrophy[12],entrophy[25],entrophy[21],datain[7]};
         20 :load =   {entrophy[24],entrophy[2],datain[0],entrophy[21],entrophy[0],entrophy[8],entrophy[11],datain[7],datain[3],datain[5],entrophy[22],entrophy[9] ,entrophy[7],entrophy[31],entrophy[15],entrophy[29],datain[2],datain[6],entrophy[12],entrophy[1],entrophy[30],entrophy[25],entrophy[23],datain[ 1],entrophy[4],entrophy[17],datain[4],entrophy[3],entrophy[20],entrophy[6],entrophy[10],entrophy[16]};
         21 :load =    { entrophy[30],datain[2],entrophy[20],entrophy[13],entrophy[28],entrophy[11],entrophy[31],entrophy[2],entrophy[0],entrophy[4],datain[7],entrophy[24] ,datain[0],datain[6],entrophy[5],datain[1],entrophy[12],datain[3],entrophy[8],entrophy[17],entrophy[9],entrophy[7],entrophy[6],datain[5],entrophy[23],entrophy[18],entrophy[16],entrophy[10],datain[4],entrophy[19],entrophy[22],entrophy[26]};
         22 :load =   {entrophy[17],entrophy[13],datain[2],entrophy[11],entrophy[16],datain[0],entrophy[3],entrophy[6],entrophy[31],entrophy[20],entrophy[7],entrophy[0] ,entrophy[27],entrophy[14],entrophy[12],entrophy[5],entrophy[21],entrophy[10],entrophy[9],datain[7],entrophy[1],entrophy[18],entrophy[22],entrophy[23],entrophy[26],datain[4],entrophy[4],datain[6],entrophy[15],datain[3],datain[1],datain[5]};
         23 :load =   {entrophy[19],datain[1],entrophy[8],entrophy[23],datain[7],datain[2],entrophy[7],datain[3],entrophy[5],entrophy[28],datain[4] ,entrophy[20],entrophy[17],entrophy[2],entrophy[16],datain[6],datain[5],entrophy[14],entrophy[30],entrophy[1],entrophy[9],datain[0],entrophy[13 ],entrophy[10],entrophy[24],entrophy[11],entrophy[0],entrophy[12],entrophy[4],entrophy[26],entrophy[3],entrophy[29]};
         24 :load =   {entrophy[16],entrophy[2],entrophy[26],entrophy[14],datain[1],entrophy[7],entrophy[1],datain[6],entrophy[18],entrophy[23],entrophy[20],datain[2] ,entrophy[30],entrophy[21],entrophy[3],entrophy[8],entrophy[31],entrophy[11],entrophy[19],entrophy[24],datain[3],entrophy[6],entrophy[4],datain[0],datain[5],entrophy[29],entrophy[12],datain[7],datain[4],entrophy[28],entrophy[17],entrophy[15] };
         25 :load =   {entrophy[31],datain[0],datain[2],entrophy[30],entrophy[9],entrophy[27],entrophy[29],entrophy[22],entrophy[13],entrophy[3],datain[6],entrophy[12] ,entrophy[0],datain[4],entrophy[19],entrophy[6],datain[7],entrophy[16],entrophy[20],entrophy[18],datain[5],entrophy[7],entrophy[10],entrophy[14 ],entrophy[25],entrophy[8],datain[1],entrophy[17],entrophy[1],entrophy[15],datain[3],entrophy[24]};
         26 :load =   {entrophy[3],entrophy[13],datain[4],entrophy[12],entrophy[14],datain[7],entrophy[0],datain[0],entrophy[20],entrophy[26],entrophy[16],datain[6] ,entrophy[19],datain[1],entrophy[11],entrophy[10],entrophy[18],datain[2],entrophy[1],entrophy[23],entrophy[7],entrophy[17],entrophy[29],entrophy[2],entrophy[27],entrophy[4],entrophy[8],datain[3],entrophy[31],entrophy[30],entrophy[5],datain[5]};
         27 :load =   {datain[2],entrophy[9],entrophy[24],entrophy[18],entrophy[23],entrophy[1],datain[0],entrophy[12],entrophy[28],entrophy[30],entrophy[17],entrophy[6] ,entrophy[5],entrophy[2],datain[3],entrophy[8],entrophy[26],datain[6],datain[4],entrophy[21],datain[1],datain[7],datain[5 ],entrophy[19],entrophy[7],entrophy[27],entrophy[0],entrophy[22],entrophy[13],entrophy[31],entrophy[15],entrophy[25]};
         28 :load =    {entrophy[26],datain[1],entrophy[9],datain[5],entrophy[2],entrophy[18],entrophy[27],datain[3],entrophy[20],entrophy[23],entrophy[4],entrophy[15] ,datain[2],entrophy[8],datain[7],datain[6],entrophy[22],entrophy[11],entrophy[6],entrophy[28],entrophy[16],entrophy[21],entrophy[7],entrophy[12 ],entrophy[14],entrophy[25],entrophy[13],entrophy[5],datain[0],entrophy[17],entrophy[0],datain[4] };
         29 :load =    {entrophy[14],entrophy[31],entrophy[18],entrophy[26],entrophy[23],entrophy[22],entrophy[24],entrophy[13],entrophy[25],datain[0],datain[6],datain[4] ,entrophy[27],entrophy[0],datain[3],entrophy[11],datain[7],datain[1],entrophy[20],entrophy[17],entrophy[29],entrophy[30],entrophy[4],entrophy[19],datain[2],entrophy[9],entrophy[2],entrophy[28],entrophy[8],entrophy[10],entrophy[7],datain[5] };
         30 :load =    {entrophy[23],datain[1],entrophy[30],datain[3],entrophy[12],entrophy[10],entrophy[6],entrophy[15],entrophy[4],entrophy[28],entrophy[5],entrophy[3] ,entrophy[14],entrophy[7],entrophy[11],entrophy[2],entrophy[17],entrophy[9],datain[0],entrophy[1],entrophy[26],datain[6],entrophy[22],entrophy[8],datain[5],datain[7],datain[2],entrophy[13],entrophy[25],entrophy[21],entrophy[16],datain[4] };
         31 :load =   {datain[0],datain[7],entrophy[8],datain[6],entrophy[14],datain[4],entrophy[24],entrophy[3],entrophy[21],entrophy[29],datain[2] ,datain[3],entrophy[0],entrophy[30],entrophy[9],datain[1],entrophy[15],entrophy[6],entrophy[17],entrophy[16],datain[5],entrophy[1],entrophy[25],entrophy[2],entrophy[11],entrophy[18],entrophy[5],entrophy[22],entrophy[4],entrophy[19],entrophy[20],entrophy[27]};
      endcase 
end    

endmodule

